magic
tech sky130A
magscale 1 2
timestamp 1699003216
<< obsli1 >>
rect 1104 2159 6532 7633
<< obsm1 >>
rect 1104 2128 6794 7664
<< metal2 >>
rect 18 0 74 800
rect 662 0 718 800
<< obsm2 >>
rect 1628 2139 6790 7653
<< metal3 >>
rect 6888 6128 7688 6248
rect 6888 5448 7688 5568
rect 6888 4768 7688 4888
rect 6888 4088 7688 4208
<< obsm3 >>
rect 1624 6328 6888 7649
rect 1624 6048 6808 6328
rect 1624 5648 6888 6048
rect 1624 5368 6808 5648
rect 1624 4968 6888 5368
rect 1624 4688 6808 4968
rect 1624 4288 6888 4688
rect 1624 4008 6808 4288
rect 1624 2143 6888 4008
<< metal4 >>
rect 1622 2128 1942 7664
rect 2282 2128 2602 7752
rect 2978 2128 3298 7664
rect 3638 2128 3958 7752
rect 4334 2128 4654 7664
rect 4994 2128 5314 7752
rect 5690 2128 6010 7664
rect 6350 2128 6670 7752
<< metal5 >>
rect 1056 7432 6670 7752
rect 1056 6772 6580 7092
rect 1056 6073 6670 6393
rect 1056 5413 6580 5733
rect 1056 4714 6670 5034
rect 1056 4054 6580 4374
rect 1056 3355 6670 3675
rect 1056 2695 6580 3015
<< labels >>
rlabel metal4 s 2282 2128 2602 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3638 2128 3958 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4994 2128 5314 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6350 2128 6670 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3355 6670 3675 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4714 6670 5034 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6073 6670 6393 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7432 6670 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1622 2128 1942 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 2978 2128 3298 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4334 2128 4654 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5690 2128 6010 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2695 6580 3015 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4054 6580 4374 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5413 6580 5733 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6772 6580 7092 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 18 0 74 800 6 b
port 3 nsew signal input
rlabel metal2 s 662 0 718 800 6 clk
port 4 nsew signal input
rlabel metal3 s 6888 6128 7688 6248 6 q[0]
port 5 nsew signal output
rlabel metal3 s 6888 4768 7688 4888 6 q[1]
port 6 nsew signal output
rlabel metal3 s 6888 4088 7688 4208 6 q[2]
port 7 nsew signal output
rlabel metal3 s 6888 5448 7688 5568 6 q[3]
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 7688 9832
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 77090
string GDS_FILE /openlane/designs/sipo/runs/RUN_2023.11.03_09.17.27/results/signoff/pes_sipo.magic.gds
string GDS_START 17080
<< end >>

