magic
tech sky130A
magscale 1 2
timestamp 1699003244
<< checkpaint >>
rect -3914 -3932 11620 11684
<< viali >>
rect 6193 6137 6227 6171
rect 6193 5661 6227 5695
rect 6193 4981 6227 5015
rect 6193 4573 6227 4607
<< metal1 >>
rect 1104 7642 6670 7664
rect 1104 7590 2288 7642
rect 2340 7590 2352 7642
rect 2404 7590 2416 7642
rect 2468 7590 2480 7642
rect 2532 7590 2544 7642
rect 2596 7590 3644 7642
rect 3696 7590 3708 7642
rect 3760 7590 3772 7642
rect 3824 7590 3836 7642
rect 3888 7590 3900 7642
rect 3952 7590 5000 7642
rect 5052 7590 5064 7642
rect 5116 7590 5128 7642
rect 5180 7590 5192 7642
rect 5244 7590 5256 7642
rect 5308 7590 6356 7642
rect 6408 7590 6420 7642
rect 6472 7590 6484 7642
rect 6536 7590 6548 7642
rect 6600 7590 6612 7642
rect 6664 7590 6670 7642
rect 1104 7568 6670 7590
rect 1104 7098 6532 7120
rect 1104 7046 1628 7098
rect 1680 7046 1692 7098
rect 1744 7046 1756 7098
rect 1808 7046 1820 7098
rect 1872 7046 1884 7098
rect 1936 7046 2984 7098
rect 3036 7046 3048 7098
rect 3100 7046 3112 7098
rect 3164 7046 3176 7098
rect 3228 7046 3240 7098
rect 3292 7046 4340 7098
rect 4392 7046 4404 7098
rect 4456 7046 4468 7098
rect 4520 7046 4532 7098
rect 4584 7046 4596 7098
rect 4648 7046 5696 7098
rect 5748 7046 5760 7098
rect 5812 7046 5824 7098
rect 5876 7046 5888 7098
rect 5940 7046 5952 7098
rect 6004 7046 6532 7098
rect 1104 7024 6532 7046
rect 1104 6554 6670 6576
rect 1104 6502 2288 6554
rect 2340 6502 2352 6554
rect 2404 6502 2416 6554
rect 2468 6502 2480 6554
rect 2532 6502 2544 6554
rect 2596 6502 3644 6554
rect 3696 6502 3708 6554
rect 3760 6502 3772 6554
rect 3824 6502 3836 6554
rect 3888 6502 3900 6554
rect 3952 6502 5000 6554
rect 5052 6502 5064 6554
rect 5116 6502 5128 6554
rect 5180 6502 5192 6554
rect 5244 6502 5256 6554
rect 5308 6502 6356 6554
rect 6408 6502 6420 6554
rect 6472 6502 6484 6554
rect 6536 6502 6548 6554
rect 6600 6502 6612 6554
rect 6664 6502 6670 6554
rect 1104 6480 6670 6502
rect 6178 6128 6184 6180
rect 6236 6128 6242 6180
rect 1104 6010 6532 6032
rect 1104 5958 1628 6010
rect 1680 5958 1692 6010
rect 1744 5958 1756 6010
rect 1808 5958 1820 6010
rect 1872 5958 1884 6010
rect 1936 5958 2984 6010
rect 3036 5958 3048 6010
rect 3100 5958 3112 6010
rect 3164 5958 3176 6010
rect 3228 5958 3240 6010
rect 3292 5958 4340 6010
rect 4392 5958 4404 6010
rect 4456 5958 4468 6010
rect 4520 5958 4532 6010
rect 4584 5958 4596 6010
rect 4648 5958 5696 6010
rect 5748 5958 5760 6010
rect 5812 5958 5824 6010
rect 5876 5958 5888 6010
rect 5940 5958 5952 6010
rect 6004 5958 6532 6010
rect 1104 5936 6532 5958
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 6730 5692 6736 5704
rect 6227 5664 6736 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 1104 5466 6670 5488
rect 1104 5414 2288 5466
rect 2340 5414 2352 5466
rect 2404 5414 2416 5466
rect 2468 5414 2480 5466
rect 2532 5414 2544 5466
rect 2596 5414 3644 5466
rect 3696 5414 3708 5466
rect 3760 5414 3772 5466
rect 3824 5414 3836 5466
rect 3888 5414 3900 5466
rect 3952 5414 5000 5466
rect 5052 5414 5064 5466
rect 5116 5414 5128 5466
rect 5180 5414 5192 5466
rect 5244 5414 5256 5466
rect 5308 5414 6356 5466
rect 6408 5414 6420 5466
rect 6472 5414 6484 5466
rect 6536 5414 6548 5466
rect 6600 5414 6612 5466
rect 6664 5414 6670 5466
rect 1104 5392 6670 5414
rect 6178 4972 6184 5024
rect 6236 4972 6242 5024
rect 1104 4922 6532 4944
rect 1104 4870 1628 4922
rect 1680 4870 1692 4922
rect 1744 4870 1756 4922
rect 1808 4870 1820 4922
rect 1872 4870 1884 4922
rect 1936 4870 2984 4922
rect 3036 4870 3048 4922
rect 3100 4870 3112 4922
rect 3164 4870 3176 4922
rect 3228 4870 3240 4922
rect 3292 4870 4340 4922
rect 4392 4870 4404 4922
rect 4456 4870 4468 4922
rect 4520 4870 4532 4922
rect 4584 4870 4596 4922
rect 4648 4870 5696 4922
rect 5748 4870 5760 4922
rect 5812 4870 5824 4922
rect 5876 4870 5888 4922
rect 5940 4870 5952 4922
rect 6004 4870 6532 4922
rect 1104 4848 6532 4870
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 1104 4378 6670 4400
rect 1104 4326 2288 4378
rect 2340 4326 2352 4378
rect 2404 4326 2416 4378
rect 2468 4326 2480 4378
rect 2532 4326 2544 4378
rect 2596 4326 3644 4378
rect 3696 4326 3708 4378
rect 3760 4326 3772 4378
rect 3824 4326 3836 4378
rect 3888 4326 3900 4378
rect 3952 4326 5000 4378
rect 5052 4326 5064 4378
rect 5116 4326 5128 4378
rect 5180 4326 5192 4378
rect 5244 4326 5256 4378
rect 5308 4326 6356 4378
rect 6408 4326 6420 4378
rect 6472 4326 6484 4378
rect 6536 4326 6548 4378
rect 6600 4326 6612 4378
rect 6664 4326 6670 4378
rect 1104 4304 6670 4326
rect 1104 3834 6532 3856
rect 1104 3782 1628 3834
rect 1680 3782 1692 3834
rect 1744 3782 1756 3834
rect 1808 3782 1820 3834
rect 1872 3782 1884 3834
rect 1936 3782 2984 3834
rect 3036 3782 3048 3834
rect 3100 3782 3112 3834
rect 3164 3782 3176 3834
rect 3228 3782 3240 3834
rect 3292 3782 4340 3834
rect 4392 3782 4404 3834
rect 4456 3782 4468 3834
rect 4520 3782 4532 3834
rect 4584 3782 4596 3834
rect 4648 3782 5696 3834
rect 5748 3782 5760 3834
rect 5812 3782 5824 3834
rect 5876 3782 5888 3834
rect 5940 3782 5952 3834
rect 6004 3782 6532 3834
rect 1104 3760 6532 3782
rect 1104 3290 6670 3312
rect 1104 3238 2288 3290
rect 2340 3238 2352 3290
rect 2404 3238 2416 3290
rect 2468 3238 2480 3290
rect 2532 3238 2544 3290
rect 2596 3238 3644 3290
rect 3696 3238 3708 3290
rect 3760 3238 3772 3290
rect 3824 3238 3836 3290
rect 3888 3238 3900 3290
rect 3952 3238 5000 3290
rect 5052 3238 5064 3290
rect 5116 3238 5128 3290
rect 5180 3238 5192 3290
rect 5244 3238 5256 3290
rect 5308 3238 6356 3290
rect 6408 3238 6420 3290
rect 6472 3238 6484 3290
rect 6536 3238 6548 3290
rect 6600 3238 6612 3290
rect 6664 3238 6670 3290
rect 1104 3216 6670 3238
rect 1104 2746 6532 2768
rect 1104 2694 1628 2746
rect 1680 2694 1692 2746
rect 1744 2694 1756 2746
rect 1808 2694 1820 2746
rect 1872 2694 1884 2746
rect 1936 2694 2984 2746
rect 3036 2694 3048 2746
rect 3100 2694 3112 2746
rect 3164 2694 3176 2746
rect 3228 2694 3240 2746
rect 3292 2694 4340 2746
rect 4392 2694 4404 2746
rect 4456 2694 4468 2746
rect 4520 2694 4532 2746
rect 4584 2694 4596 2746
rect 4648 2694 5696 2746
rect 5748 2694 5760 2746
rect 5812 2694 5824 2746
rect 5876 2694 5888 2746
rect 5940 2694 5952 2746
rect 6004 2694 6532 2746
rect 1104 2672 6532 2694
rect 1104 2202 6670 2224
rect 1104 2150 2288 2202
rect 2340 2150 2352 2202
rect 2404 2150 2416 2202
rect 2468 2150 2480 2202
rect 2532 2150 2544 2202
rect 2596 2150 3644 2202
rect 3696 2150 3708 2202
rect 3760 2150 3772 2202
rect 3824 2150 3836 2202
rect 3888 2150 3900 2202
rect 3952 2150 5000 2202
rect 5052 2150 5064 2202
rect 5116 2150 5128 2202
rect 5180 2150 5192 2202
rect 5244 2150 5256 2202
rect 5308 2150 6356 2202
rect 6408 2150 6420 2202
rect 6472 2150 6484 2202
rect 6536 2150 6548 2202
rect 6600 2150 6612 2202
rect 6664 2150 6670 2202
rect 1104 2128 6670 2150
<< via1 >>
rect 2288 7590 2340 7642
rect 2352 7590 2404 7642
rect 2416 7590 2468 7642
rect 2480 7590 2532 7642
rect 2544 7590 2596 7642
rect 3644 7590 3696 7642
rect 3708 7590 3760 7642
rect 3772 7590 3824 7642
rect 3836 7590 3888 7642
rect 3900 7590 3952 7642
rect 5000 7590 5052 7642
rect 5064 7590 5116 7642
rect 5128 7590 5180 7642
rect 5192 7590 5244 7642
rect 5256 7590 5308 7642
rect 6356 7590 6408 7642
rect 6420 7590 6472 7642
rect 6484 7590 6536 7642
rect 6548 7590 6600 7642
rect 6612 7590 6664 7642
rect 1628 7046 1680 7098
rect 1692 7046 1744 7098
rect 1756 7046 1808 7098
rect 1820 7046 1872 7098
rect 1884 7046 1936 7098
rect 2984 7046 3036 7098
rect 3048 7046 3100 7098
rect 3112 7046 3164 7098
rect 3176 7046 3228 7098
rect 3240 7046 3292 7098
rect 4340 7046 4392 7098
rect 4404 7046 4456 7098
rect 4468 7046 4520 7098
rect 4532 7046 4584 7098
rect 4596 7046 4648 7098
rect 5696 7046 5748 7098
rect 5760 7046 5812 7098
rect 5824 7046 5876 7098
rect 5888 7046 5940 7098
rect 5952 7046 6004 7098
rect 2288 6502 2340 6554
rect 2352 6502 2404 6554
rect 2416 6502 2468 6554
rect 2480 6502 2532 6554
rect 2544 6502 2596 6554
rect 3644 6502 3696 6554
rect 3708 6502 3760 6554
rect 3772 6502 3824 6554
rect 3836 6502 3888 6554
rect 3900 6502 3952 6554
rect 5000 6502 5052 6554
rect 5064 6502 5116 6554
rect 5128 6502 5180 6554
rect 5192 6502 5244 6554
rect 5256 6502 5308 6554
rect 6356 6502 6408 6554
rect 6420 6502 6472 6554
rect 6484 6502 6536 6554
rect 6548 6502 6600 6554
rect 6612 6502 6664 6554
rect 6184 6171 6236 6180
rect 6184 6137 6193 6171
rect 6193 6137 6227 6171
rect 6227 6137 6236 6171
rect 6184 6128 6236 6137
rect 1628 5958 1680 6010
rect 1692 5958 1744 6010
rect 1756 5958 1808 6010
rect 1820 5958 1872 6010
rect 1884 5958 1936 6010
rect 2984 5958 3036 6010
rect 3048 5958 3100 6010
rect 3112 5958 3164 6010
rect 3176 5958 3228 6010
rect 3240 5958 3292 6010
rect 4340 5958 4392 6010
rect 4404 5958 4456 6010
rect 4468 5958 4520 6010
rect 4532 5958 4584 6010
rect 4596 5958 4648 6010
rect 5696 5958 5748 6010
rect 5760 5958 5812 6010
rect 5824 5958 5876 6010
rect 5888 5958 5940 6010
rect 5952 5958 6004 6010
rect 6736 5652 6788 5704
rect 2288 5414 2340 5466
rect 2352 5414 2404 5466
rect 2416 5414 2468 5466
rect 2480 5414 2532 5466
rect 2544 5414 2596 5466
rect 3644 5414 3696 5466
rect 3708 5414 3760 5466
rect 3772 5414 3824 5466
rect 3836 5414 3888 5466
rect 3900 5414 3952 5466
rect 5000 5414 5052 5466
rect 5064 5414 5116 5466
rect 5128 5414 5180 5466
rect 5192 5414 5244 5466
rect 5256 5414 5308 5466
rect 6356 5414 6408 5466
rect 6420 5414 6472 5466
rect 6484 5414 6536 5466
rect 6548 5414 6600 5466
rect 6612 5414 6664 5466
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 1628 4870 1680 4922
rect 1692 4870 1744 4922
rect 1756 4870 1808 4922
rect 1820 4870 1872 4922
rect 1884 4870 1936 4922
rect 2984 4870 3036 4922
rect 3048 4870 3100 4922
rect 3112 4870 3164 4922
rect 3176 4870 3228 4922
rect 3240 4870 3292 4922
rect 4340 4870 4392 4922
rect 4404 4870 4456 4922
rect 4468 4870 4520 4922
rect 4532 4870 4584 4922
rect 4596 4870 4648 4922
rect 5696 4870 5748 4922
rect 5760 4870 5812 4922
rect 5824 4870 5876 4922
rect 5888 4870 5940 4922
rect 5952 4870 6004 4922
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 2288 4326 2340 4378
rect 2352 4326 2404 4378
rect 2416 4326 2468 4378
rect 2480 4326 2532 4378
rect 2544 4326 2596 4378
rect 3644 4326 3696 4378
rect 3708 4326 3760 4378
rect 3772 4326 3824 4378
rect 3836 4326 3888 4378
rect 3900 4326 3952 4378
rect 5000 4326 5052 4378
rect 5064 4326 5116 4378
rect 5128 4326 5180 4378
rect 5192 4326 5244 4378
rect 5256 4326 5308 4378
rect 6356 4326 6408 4378
rect 6420 4326 6472 4378
rect 6484 4326 6536 4378
rect 6548 4326 6600 4378
rect 6612 4326 6664 4378
rect 1628 3782 1680 3834
rect 1692 3782 1744 3834
rect 1756 3782 1808 3834
rect 1820 3782 1872 3834
rect 1884 3782 1936 3834
rect 2984 3782 3036 3834
rect 3048 3782 3100 3834
rect 3112 3782 3164 3834
rect 3176 3782 3228 3834
rect 3240 3782 3292 3834
rect 4340 3782 4392 3834
rect 4404 3782 4456 3834
rect 4468 3782 4520 3834
rect 4532 3782 4584 3834
rect 4596 3782 4648 3834
rect 5696 3782 5748 3834
rect 5760 3782 5812 3834
rect 5824 3782 5876 3834
rect 5888 3782 5940 3834
rect 5952 3782 6004 3834
rect 2288 3238 2340 3290
rect 2352 3238 2404 3290
rect 2416 3238 2468 3290
rect 2480 3238 2532 3290
rect 2544 3238 2596 3290
rect 3644 3238 3696 3290
rect 3708 3238 3760 3290
rect 3772 3238 3824 3290
rect 3836 3238 3888 3290
rect 3900 3238 3952 3290
rect 5000 3238 5052 3290
rect 5064 3238 5116 3290
rect 5128 3238 5180 3290
rect 5192 3238 5244 3290
rect 5256 3238 5308 3290
rect 6356 3238 6408 3290
rect 6420 3238 6472 3290
rect 6484 3238 6536 3290
rect 6548 3238 6600 3290
rect 6612 3238 6664 3290
rect 1628 2694 1680 2746
rect 1692 2694 1744 2746
rect 1756 2694 1808 2746
rect 1820 2694 1872 2746
rect 1884 2694 1936 2746
rect 2984 2694 3036 2746
rect 3048 2694 3100 2746
rect 3112 2694 3164 2746
rect 3176 2694 3228 2746
rect 3240 2694 3292 2746
rect 4340 2694 4392 2746
rect 4404 2694 4456 2746
rect 4468 2694 4520 2746
rect 4532 2694 4584 2746
rect 4596 2694 4648 2746
rect 5696 2694 5748 2746
rect 5760 2694 5812 2746
rect 5824 2694 5876 2746
rect 5888 2694 5940 2746
rect 5952 2694 6004 2746
rect 2288 2150 2340 2202
rect 2352 2150 2404 2202
rect 2416 2150 2468 2202
rect 2480 2150 2532 2202
rect 2544 2150 2596 2202
rect 3644 2150 3696 2202
rect 3708 2150 3760 2202
rect 3772 2150 3824 2202
rect 3836 2150 3888 2202
rect 3900 2150 3952 2202
rect 5000 2150 5052 2202
rect 5064 2150 5116 2202
rect 5128 2150 5180 2202
rect 5192 2150 5244 2202
rect 5256 2150 5308 2202
rect 6356 2150 6408 2202
rect 6420 2150 6472 2202
rect 6484 2150 6536 2202
rect 6548 2150 6600 2202
rect 6612 2150 6664 2202
<< metal2 >>
rect 2288 7644 2596 7653
rect 2288 7642 2294 7644
rect 2350 7642 2374 7644
rect 2430 7642 2454 7644
rect 2510 7642 2534 7644
rect 2590 7642 2596 7644
rect 2350 7590 2352 7642
rect 2532 7590 2534 7642
rect 2288 7588 2294 7590
rect 2350 7588 2374 7590
rect 2430 7588 2454 7590
rect 2510 7588 2534 7590
rect 2590 7588 2596 7590
rect 2288 7579 2596 7588
rect 3644 7644 3952 7653
rect 3644 7642 3650 7644
rect 3706 7642 3730 7644
rect 3786 7642 3810 7644
rect 3866 7642 3890 7644
rect 3946 7642 3952 7644
rect 3706 7590 3708 7642
rect 3888 7590 3890 7642
rect 3644 7588 3650 7590
rect 3706 7588 3730 7590
rect 3786 7588 3810 7590
rect 3866 7588 3890 7590
rect 3946 7588 3952 7590
rect 3644 7579 3952 7588
rect 5000 7644 5308 7653
rect 5000 7642 5006 7644
rect 5062 7642 5086 7644
rect 5142 7642 5166 7644
rect 5222 7642 5246 7644
rect 5302 7642 5308 7644
rect 5062 7590 5064 7642
rect 5244 7590 5246 7642
rect 5000 7588 5006 7590
rect 5062 7588 5086 7590
rect 5142 7588 5166 7590
rect 5222 7588 5246 7590
rect 5302 7588 5308 7590
rect 5000 7579 5308 7588
rect 6356 7644 6664 7653
rect 6356 7642 6362 7644
rect 6418 7642 6442 7644
rect 6498 7642 6522 7644
rect 6578 7642 6602 7644
rect 6658 7642 6664 7644
rect 6418 7590 6420 7642
rect 6600 7590 6602 7642
rect 6356 7588 6362 7590
rect 6418 7588 6442 7590
rect 6498 7588 6522 7590
rect 6578 7588 6602 7590
rect 6658 7588 6664 7590
rect 6356 7579 6664 7588
rect 1628 7100 1936 7109
rect 1628 7098 1634 7100
rect 1690 7098 1714 7100
rect 1770 7098 1794 7100
rect 1850 7098 1874 7100
rect 1930 7098 1936 7100
rect 1690 7046 1692 7098
rect 1872 7046 1874 7098
rect 1628 7044 1634 7046
rect 1690 7044 1714 7046
rect 1770 7044 1794 7046
rect 1850 7044 1874 7046
rect 1930 7044 1936 7046
rect 1628 7035 1936 7044
rect 2984 7100 3292 7109
rect 2984 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3150 7100
rect 3206 7098 3230 7100
rect 3286 7098 3292 7100
rect 3046 7046 3048 7098
rect 3228 7046 3230 7098
rect 2984 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3150 7046
rect 3206 7044 3230 7046
rect 3286 7044 3292 7046
rect 2984 7035 3292 7044
rect 4340 7100 4648 7109
rect 4340 7098 4346 7100
rect 4402 7098 4426 7100
rect 4482 7098 4506 7100
rect 4562 7098 4586 7100
rect 4642 7098 4648 7100
rect 4402 7046 4404 7098
rect 4584 7046 4586 7098
rect 4340 7044 4346 7046
rect 4402 7044 4426 7046
rect 4482 7044 4506 7046
rect 4562 7044 4586 7046
rect 4642 7044 4648 7046
rect 4340 7035 4648 7044
rect 5696 7100 6004 7109
rect 5696 7098 5702 7100
rect 5758 7098 5782 7100
rect 5838 7098 5862 7100
rect 5918 7098 5942 7100
rect 5998 7098 6004 7100
rect 5758 7046 5760 7098
rect 5940 7046 5942 7098
rect 5696 7044 5702 7046
rect 5758 7044 5782 7046
rect 5838 7044 5862 7046
rect 5918 7044 5942 7046
rect 5998 7044 6004 7046
rect 5696 7035 6004 7044
rect 2288 6556 2596 6565
rect 2288 6554 2294 6556
rect 2350 6554 2374 6556
rect 2430 6554 2454 6556
rect 2510 6554 2534 6556
rect 2590 6554 2596 6556
rect 2350 6502 2352 6554
rect 2532 6502 2534 6554
rect 2288 6500 2294 6502
rect 2350 6500 2374 6502
rect 2430 6500 2454 6502
rect 2510 6500 2534 6502
rect 2590 6500 2596 6502
rect 2288 6491 2596 6500
rect 3644 6556 3952 6565
rect 3644 6554 3650 6556
rect 3706 6554 3730 6556
rect 3786 6554 3810 6556
rect 3866 6554 3890 6556
rect 3946 6554 3952 6556
rect 3706 6502 3708 6554
rect 3888 6502 3890 6554
rect 3644 6500 3650 6502
rect 3706 6500 3730 6502
rect 3786 6500 3810 6502
rect 3866 6500 3890 6502
rect 3946 6500 3952 6502
rect 3644 6491 3952 6500
rect 5000 6556 5308 6565
rect 5000 6554 5006 6556
rect 5062 6554 5086 6556
rect 5142 6554 5166 6556
rect 5222 6554 5246 6556
rect 5302 6554 5308 6556
rect 5062 6502 5064 6554
rect 5244 6502 5246 6554
rect 5000 6500 5006 6502
rect 5062 6500 5086 6502
rect 5142 6500 5166 6502
rect 5222 6500 5246 6502
rect 5302 6500 5308 6502
rect 5000 6491 5308 6500
rect 6356 6556 6664 6565
rect 6356 6554 6362 6556
rect 6418 6554 6442 6556
rect 6498 6554 6522 6556
rect 6578 6554 6602 6556
rect 6658 6554 6664 6556
rect 6418 6502 6420 6554
rect 6600 6502 6602 6554
rect 6356 6500 6362 6502
rect 6418 6500 6442 6502
rect 6498 6500 6522 6502
rect 6578 6500 6602 6502
rect 6658 6500 6664 6502
rect 6356 6491 6664 6500
rect 6182 6216 6238 6225
rect 6182 6151 6184 6160
rect 6236 6151 6238 6160
rect 6184 6122 6236 6128
rect 1628 6012 1936 6021
rect 1628 6010 1634 6012
rect 1690 6010 1714 6012
rect 1770 6010 1794 6012
rect 1850 6010 1874 6012
rect 1930 6010 1936 6012
rect 1690 5958 1692 6010
rect 1872 5958 1874 6010
rect 1628 5956 1634 5958
rect 1690 5956 1714 5958
rect 1770 5956 1794 5958
rect 1850 5956 1874 5958
rect 1930 5956 1936 5958
rect 1628 5947 1936 5956
rect 2984 6012 3292 6021
rect 2984 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3150 6012
rect 3206 6010 3230 6012
rect 3286 6010 3292 6012
rect 3046 5958 3048 6010
rect 3228 5958 3230 6010
rect 2984 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3150 5958
rect 3206 5956 3230 5958
rect 3286 5956 3292 5958
rect 2984 5947 3292 5956
rect 4340 6012 4648 6021
rect 4340 6010 4346 6012
rect 4402 6010 4426 6012
rect 4482 6010 4506 6012
rect 4562 6010 4586 6012
rect 4642 6010 4648 6012
rect 4402 5958 4404 6010
rect 4584 5958 4586 6010
rect 4340 5956 4346 5958
rect 4402 5956 4426 5958
rect 4482 5956 4506 5958
rect 4562 5956 4586 5958
rect 4642 5956 4648 5958
rect 4340 5947 4648 5956
rect 5696 6012 6004 6021
rect 5696 6010 5702 6012
rect 5758 6010 5782 6012
rect 5838 6010 5862 6012
rect 5918 6010 5942 6012
rect 5998 6010 6004 6012
rect 5758 5958 5760 6010
rect 5940 5958 5942 6010
rect 5696 5956 5702 5958
rect 5758 5956 5782 5958
rect 5838 5956 5862 5958
rect 5918 5956 5942 5958
rect 5998 5956 6004 5958
rect 5696 5947 6004 5956
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 5545 6776 5646
rect 6734 5536 6790 5545
rect 2288 5468 2596 5477
rect 2288 5466 2294 5468
rect 2350 5466 2374 5468
rect 2430 5466 2454 5468
rect 2510 5466 2534 5468
rect 2590 5466 2596 5468
rect 2350 5414 2352 5466
rect 2532 5414 2534 5466
rect 2288 5412 2294 5414
rect 2350 5412 2374 5414
rect 2430 5412 2454 5414
rect 2510 5412 2534 5414
rect 2590 5412 2596 5414
rect 2288 5403 2596 5412
rect 3644 5468 3952 5477
rect 3644 5466 3650 5468
rect 3706 5466 3730 5468
rect 3786 5466 3810 5468
rect 3866 5466 3890 5468
rect 3946 5466 3952 5468
rect 3706 5414 3708 5466
rect 3888 5414 3890 5466
rect 3644 5412 3650 5414
rect 3706 5412 3730 5414
rect 3786 5412 3810 5414
rect 3866 5412 3890 5414
rect 3946 5412 3952 5414
rect 3644 5403 3952 5412
rect 5000 5468 5308 5477
rect 5000 5466 5006 5468
rect 5062 5466 5086 5468
rect 5142 5466 5166 5468
rect 5222 5466 5246 5468
rect 5302 5466 5308 5468
rect 5062 5414 5064 5466
rect 5244 5414 5246 5466
rect 5000 5412 5006 5414
rect 5062 5412 5086 5414
rect 5142 5412 5166 5414
rect 5222 5412 5246 5414
rect 5302 5412 5308 5414
rect 5000 5403 5308 5412
rect 6356 5468 6664 5477
rect 6734 5471 6790 5480
rect 6356 5466 6362 5468
rect 6418 5466 6442 5468
rect 6498 5466 6522 5468
rect 6578 5466 6602 5468
rect 6658 5466 6664 5468
rect 6418 5414 6420 5466
rect 6600 5414 6602 5466
rect 6356 5412 6362 5414
rect 6418 5412 6442 5414
rect 6498 5412 6522 5414
rect 6578 5412 6602 5414
rect 6658 5412 6664 5414
rect 6356 5403 6664 5412
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 1628 4924 1936 4933
rect 1628 4922 1634 4924
rect 1690 4922 1714 4924
rect 1770 4922 1794 4924
rect 1850 4922 1874 4924
rect 1930 4922 1936 4924
rect 1690 4870 1692 4922
rect 1872 4870 1874 4922
rect 1628 4868 1634 4870
rect 1690 4868 1714 4870
rect 1770 4868 1794 4870
rect 1850 4868 1874 4870
rect 1930 4868 1936 4870
rect 1628 4859 1936 4868
rect 2984 4924 3292 4933
rect 2984 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3150 4924
rect 3206 4922 3230 4924
rect 3286 4922 3292 4924
rect 3046 4870 3048 4922
rect 3228 4870 3230 4922
rect 2984 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3150 4870
rect 3206 4868 3230 4870
rect 3286 4868 3292 4870
rect 2984 4859 3292 4868
rect 4340 4924 4648 4933
rect 4340 4922 4346 4924
rect 4402 4922 4426 4924
rect 4482 4922 4506 4924
rect 4562 4922 4586 4924
rect 4642 4922 4648 4924
rect 4402 4870 4404 4922
rect 4584 4870 4586 4922
rect 4340 4868 4346 4870
rect 4402 4868 4426 4870
rect 4482 4868 4506 4870
rect 4562 4868 4586 4870
rect 4642 4868 4648 4870
rect 4340 4859 4648 4868
rect 5696 4924 6004 4933
rect 5696 4922 5702 4924
rect 5758 4922 5782 4924
rect 5838 4922 5862 4924
rect 5918 4922 5942 4924
rect 5998 4922 6004 4924
rect 5758 4870 5760 4922
rect 5940 4870 5942 4922
rect 5696 4868 5702 4870
rect 5758 4868 5782 4870
rect 5838 4868 5862 4870
rect 5918 4868 5942 4870
rect 5998 4868 6004 4870
rect 5696 4859 6004 4868
rect 6196 4865 6224 4966
rect 6182 4856 6238 4865
rect 6182 4791 6238 4800
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 2288 4380 2596 4389
rect 2288 4378 2294 4380
rect 2350 4378 2374 4380
rect 2430 4378 2454 4380
rect 2510 4378 2534 4380
rect 2590 4378 2596 4380
rect 2350 4326 2352 4378
rect 2532 4326 2534 4378
rect 2288 4324 2294 4326
rect 2350 4324 2374 4326
rect 2430 4324 2454 4326
rect 2510 4324 2534 4326
rect 2590 4324 2596 4326
rect 2288 4315 2596 4324
rect 3644 4380 3952 4389
rect 3644 4378 3650 4380
rect 3706 4378 3730 4380
rect 3786 4378 3810 4380
rect 3866 4378 3890 4380
rect 3946 4378 3952 4380
rect 3706 4326 3708 4378
rect 3888 4326 3890 4378
rect 3644 4324 3650 4326
rect 3706 4324 3730 4326
rect 3786 4324 3810 4326
rect 3866 4324 3890 4326
rect 3946 4324 3952 4326
rect 3644 4315 3952 4324
rect 5000 4380 5308 4389
rect 5000 4378 5006 4380
rect 5062 4378 5086 4380
rect 5142 4378 5166 4380
rect 5222 4378 5246 4380
rect 5302 4378 5308 4380
rect 5062 4326 5064 4378
rect 5244 4326 5246 4378
rect 5000 4324 5006 4326
rect 5062 4324 5086 4326
rect 5142 4324 5166 4326
rect 5222 4324 5246 4326
rect 5302 4324 5308 4326
rect 5000 4315 5308 4324
rect 6196 4185 6224 4558
rect 6356 4380 6664 4389
rect 6356 4378 6362 4380
rect 6418 4378 6442 4380
rect 6498 4378 6522 4380
rect 6578 4378 6602 4380
rect 6658 4378 6664 4380
rect 6418 4326 6420 4378
rect 6600 4326 6602 4378
rect 6356 4324 6362 4326
rect 6418 4324 6442 4326
rect 6498 4324 6522 4326
rect 6578 4324 6602 4326
rect 6658 4324 6664 4326
rect 6356 4315 6664 4324
rect 6182 4176 6238 4185
rect 6182 4111 6238 4120
rect 1628 3836 1936 3845
rect 1628 3834 1634 3836
rect 1690 3834 1714 3836
rect 1770 3834 1794 3836
rect 1850 3834 1874 3836
rect 1930 3834 1936 3836
rect 1690 3782 1692 3834
rect 1872 3782 1874 3834
rect 1628 3780 1634 3782
rect 1690 3780 1714 3782
rect 1770 3780 1794 3782
rect 1850 3780 1874 3782
rect 1930 3780 1936 3782
rect 1628 3771 1936 3780
rect 2984 3836 3292 3845
rect 2984 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3150 3836
rect 3206 3834 3230 3836
rect 3286 3834 3292 3836
rect 3046 3782 3048 3834
rect 3228 3782 3230 3834
rect 2984 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3150 3782
rect 3206 3780 3230 3782
rect 3286 3780 3292 3782
rect 2984 3771 3292 3780
rect 4340 3836 4648 3845
rect 4340 3834 4346 3836
rect 4402 3834 4426 3836
rect 4482 3834 4506 3836
rect 4562 3834 4586 3836
rect 4642 3834 4648 3836
rect 4402 3782 4404 3834
rect 4584 3782 4586 3834
rect 4340 3780 4346 3782
rect 4402 3780 4426 3782
rect 4482 3780 4506 3782
rect 4562 3780 4586 3782
rect 4642 3780 4648 3782
rect 4340 3771 4648 3780
rect 5696 3836 6004 3845
rect 5696 3834 5702 3836
rect 5758 3834 5782 3836
rect 5838 3834 5862 3836
rect 5918 3834 5942 3836
rect 5998 3834 6004 3836
rect 5758 3782 5760 3834
rect 5940 3782 5942 3834
rect 5696 3780 5702 3782
rect 5758 3780 5782 3782
rect 5838 3780 5862 3782
rect 5918 3780 5942 3782
rect 5998 3780 6004 3782
rect 5696 3771 6004 3780
rect 2288 3292 2596 3301
rect 2288 3290 2294 3292
rect 2350 3290 2374 3292
rect 2430 3290 2454 3292
rect 2510 3290 2534 3292
rect 2590 3290 2596 3292
rect 2350 3238 2352 3290
rect 2532 3238 2534 3290
rect 2288 3236 2294 3238
rect 2350 3236 2374 3238
rect 2430 3236 2454 3238
rect 2510 3236 2534 3238
rect 2590 3236 2596 3238
rect 2288 3227 2596 3236
rect 3644 3292 3952 3301
rect 3644 3290 3650 3292
rect 3706 3290 3730 3292
rect 3786 3290 3810 3292
rect 3866 3290 3890 3292
rect 3946 3290 3952 3292
rect 3706 3238 3708 3290
rect 3888 3238 3890 3290
rect 3644 3236 3650 3238
rect 3706 3236 3730 3238
rect 3786 3236 3810 3238
rect 3866 3236 3890 3238
rect 3946 3236 3952 3238
rect 3644 3227 3952 3236
rect 5000 3292 5308 3301
rect 5000 3290 5006 3292
rect 5062 3290 5086 3292
rect 5142 3290 5166 3292
rect 5222 3290 5246 3292
rect 5302 3290 5308 3292
rect 5062 3238 5064 3290
rect 5244 3238 5246 3290
rect 5000 3236 5006 3238
rect 5062 3236 5086 3238
rect 5142 3236 5166 3238
rect 5222 3236 5246 3238
rect 5302 3236 5308 3238
rect 5000 3227 5308 3236
rect 6356 3292 6664 3301
rect 6356 3290 6362 3292
rect 6418 3290 6442 3292
rect 6498 3290 6522 3292
rect 6578 3290 6602 3292
rect 6658 3290 6664 3292
rect 6418 3238 6420 3290
rect 6600 3238 6602 3290
rect 6356 3236 6362 3238
rect 6418 3236 6442 3238
rect 6498 3236 6522 3238
rect 6578 3236 6602 3238
rect 6658 3236 6664 3238
rect 6356 3227 6664 3236
rect 1628 2748 1936 2757
rect 1628 2746 1634 2748
rect 1690 2746 1714 2748
rect 1770 2746 1794 2748
rect 1850 2746 1874 2748
rect 1930 2746 1936 2748
rect 1690 2694 1692 2746
rect 1872 2694 1874 2746
rect 1628 2692 1634 2694
rect 1690 2692 1714 2694
rect 1770 2692 1794 2694
rect 1850 2692 1874 2694
rect 1930 2692 1936 2694
rect 1628 2683 1936 2692
rect 2984 2748 3292 2757
rect 2984 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3150 2748
rect 3206 2746 3230 2748
rect 3286 2746 3292 2748
rect 3046 2694 3048 2746
rect 3228 2694 3230 2746
rect 2984 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3150 2694
rect 3206 2692 3230 2694
rect 3286 2692 3292 2694
rect 2984 2683 3292 2692
rect 4340 2748 4648 2757
rect 4340 2746 4346 2748
rect 4402 2746 4426 2748
rect 4482 2746 4506 2748
rect 4562 2746 4586 2748
rect 4642 2746 4648 2748
rect 4402 2694 4404 2746
rect 4584 2694 4586 2746
rect 4340 2692 4346 2694
rect 4402 2692 4426 2694
rect 4482 2692 4506 2694
rect 4562 2692 4586 2694
rect 4642 2692 4648 2694
rect 4340 2683 4648 2692
rect 5696 2748 6004 2757
rect 5696 2746 5702 2748
rect 5758 2746 5782 2748
rect 5838 2746 5862 2748
rect 5918 2746 5942 2748
rect 5998 2746 6004 2748
rect 5758 2694 5760 2746
rect 5940 2694 5942 2746
rect 5696 2692 5702 2694
rect 5758 2692 5782 2694
rect 5838 2692 5862 2694
rect 5918 2692 5942 2694
rect 5998 2692 6004 2694
rect 5696 2683 6004 2692
rect 2288 2204 2596 2213
rect 2288 2202 2294 2204
rect 2350 2202 2374 2204
rect 2430 2202 2454 2204
rect 2510 2202 2534 2204
rect 2590 2202 2596 2204
rect 2350 2150 2352 2202
rect 2532 2150 2534 2202
rect 2288 2148 2294 2150
rect 2350 2148 2374 2150
rect 2430 2148 2454 2150
rect 2510 2148 2534 2150
rect 2590 2148 2596 2150
rect 2288 2139 2596 2148
rect 3644 2204 3952 2213
rect 3644 2202 3650 2204
rect 3706 2202 3730 2204
rect 3786 2202 3810 2204
rect 3866 2202 3890 2204
rect 3946 2202 3952 2204
rect 3706 2150 3708 2202
rect 3888 2150 3890 2202
rect 3644 2148 3650 2150
rect 3706 2148 3730 2150
rect 3786 2148 3810 2150
rect 3866 2148 3890 2150
rect 3946 2148 3952 2150
rect 3644 2139 3952 2148
rect 5000 2204 5308 2213
rect 5000 2202 5006 2204
rect 5062 2202 5086 2204
rect 5142 2202 5166 2204
rect 5222 2202 5246 2204
rect 5302 2202 5308 2204
rect 5062 2150 5064 2202
rect 5244 2150 5246 2202
rect 5000 2148 5006 2150
rect 5062 2148 5086 2150
rect 5142 2148 5166 2150
rect 5222 2148 5246 2150
rect 5302 2148 5308 2150
rect 5000 2139 5308 2148
rect 6356 2204 6664 2213
rect 6356 2202 6362 2204
rect 6418 2202 6442 2204
rect 6498 2202 6522 2204
rect 6578 2202 6602 2204
rect 6658 2202 6664 2204
rect 6418 2150 6420 2202
rect 6600 2150 6602 2202
rect 6356 2148 6362 2150
rect 6418 2148 6442 2150
rect 6498 2148 6522 2150
rect 6578 2148 6602 2150
rect 6658 2148 6664 2150
rect 6356 2139 6664 2148
rect 18 0 74 800
rect 662 0 718 800
<< via2 >>
rect 2294 7642 2350 7644
rect 2374 7642 2430 7644
rect 2454 7642 2510 7644
rect 2534 7642 2590 7644
rect 2294 7590 2340 7642
rect 2340 7590 2350 7642
rect 2374 7590 2404 7642
rect 2404 7590 2416 7642
rect 2416 7590 2430 7642
rect 2454 7590 2468 7642
rect 2468 7590 2480 7642
rect 2480 7590 2510 7642
rect 2534 7590 2544 7642
rect 2544 7590 2590 7642
rect 2294 7588 2350 7590
rect 2374 7588 2430 7590
rect 2454 7588 2510 7590
rect 2534 7588 2590 7590
rect 3650 7642 3706 7644
rect 3730 7642 3786 7644
rect 3810 7642 3866 7644
rect 3890 7642 3946 7644
rect 3650 7590 3696 7642
rect 3696 7590 3706 7642
rect 3730 7590 3760 7642
rect 3760 7590 3772 7642
rect 3772 7590 3786 7642
rect 3810 7590 3824 7642
rect 3824 7590 3836 7642
rect 3836 7590 3866 7642
rect 3890 7590 3900 7642
rect 3900 7590 3946 7642
rect 3650 7588 3706 7590
rect 3730 7588 3786 7590
rect 3810 7588 3866 7590
rect 3890 7588 3946 7590
rect 5006 7642 5062 7644
rect 5086 7642 5142 7644
rect 5166 7642 5222 7644
rect 5246 7642 5302 7644
rect 5006 7590 5052 7642
rect 5052 7590 5062 7642
rect 5086 7590 5116 7642
rect 5116 7590 5128 7642
rect 5128 7590 5142 7642
rect 5166 7590 5180 7642
rect 5180 7590 5192 7642
rect 5192 7590 5222 7642
rect 5246 7590 5256 7642
rect 5256 7590 5302 7642
rect 5006 7588 5062 7590
rect 5086 7588 5142 7590
rect 5166 7588 5222 7590
rect 5246 7588 5302 7590
rect 6362 7642 6418 7644
rect 6442 7642 6498 7644
rect 6522 7642 6578 7644
rect 6602 7642 6658 7644
rect 6362 7590 6408 7642
rect 6408 7590 6418 7642
rect 6442 7590 6472 7642
rect 6472 7590 6484 7642
rect 6484 7590 6498 7642
rect 6522 7590 6536 7642
rect 6536 7590 6548 7642
rect 6548 7590 6578 7642
rect 6602 7590 6612 7642
rect 6612 7590 6658 7642
rect 6362 7588 6418 7590
rect 6442 7588 6498 7590
rect 6522 7588 6578 7590
rect 6602 7588 6658 7590
rect 1634 7098 1690 7100
rect 1714 7098 1770 7100
rect 1794 7098 1850 7100
rect 1874 7098 1930 7100
rect 1634 7046 1680 7098
rect 1680 7046 1690 7098
rect 1714 7046 1744 7098
rect 1744 7046 1756 7098
rect 1756 7046 1770 7098
rect 1794 7046 1808 7098
rect 1808 7046 1820 7098
rect 1820 7046 1850 7098
rect 1874 7046 1884 7098
rect 1884 7046 1930 7098
rect 1634 7044 1690 7046
rect 1714 7044 1770 7046
rect 1794 7044 1850 7046
rect 1874 7044 1930 7046
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 3150 7098 3206 7100
rect 3230 7098 3286 7100
rect 2990 7046 3036 7098
rect 3036 7046 3046 7098
rect 3070 7046 3100 7098
rect 3100 7046 3112 7098
rect 3112 7046 3126 7098
rect 3150 7046 3164 7098
rect 3164 7046 3176 7098
rect 3176 7046 3206 7098
rect 3230 7046 3240 7098
rect 3240 7046 3286 7098
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 3150 7044 3206 7046
rect 3230 7044 3286 7046
rect 4346 7098 4402 7100
rect 4426 7098 4482 7100
rect 4506 7098 4562 7100
rect 4586 7098 4642 7100
rect 4346 7046 4392 7098
rect 4392 7046 4402 7098
rect 4426 7046 4456 7098
rect 4456 7046 4468 7098
rect 4468 7046 4482 7098
rect 4506 7046 4520 7098
rect 4520 7046 4532 7098
rect 4532 7046 4562 7098
rect 4586 7046 4596 7098
rect 4596 7046 4642 7098
rect 4346 7044 4402 7046
rect 4426 7044 4482 7046
rect 4506 7044 4562 7046
rect 4586 7044 4642 7046
rect 5702 7098 5758 7100
rect 5782 7098 5838 7100
rect 5862 7098 5918 7100
rect 5942 7098 5998 7100
rect 5702 7046 5748 7098
rect 5748 7046 5758 7098
rect 5782 7046 5812 7098
rect 5812 7046 5824 7098
rect 5824 7046 5838 7098
rect 5862 7046 5876 7098
rect 5876 7046 5888 7098
rect 5888 7046 5918 7098
rect 5942 7046 5952 7098
rect 5952 7046 5998 7098
rect 5702 7044 5758 7046
rect 5782 7044 5838 7046
rect 5862 7044 5918 7046
rect 5942 7044 5998 7046
rect 2294 6554 2350 6556
rect 2374 6554 2430 6556
rect 2454 6554 2510 6556
rect 2534 6554 2590 6556
rect 2294 6502 2340 6554
rect 2340 6502 2350 6554
rect 2374 6502 2404 6554
rect 2404 6502 2416 6554
rect 2416 6502 2430 6554
rect 2454 6502 2468 6554
rect 2468 6502 2480 6554
rect 2480 6502 2510 6554
rect 2534 6502 2544 6554
rect 2544 6502 2590 6554
rect 2294 6500 2350 6502
rect 2374 6500 2430 6502
rect 2454 6500 2510 6502
rect 2534 6500 2590 6502
rect 3650 6554 3706 6556
rect 3730 6554 3786 6556
rect 3810 6554 3866 6556
rect 3890 6554 3946 6556
rect 3650 6502 3696 6554
rect 3696 6502 3706 6554
rect 3730 6502 3760 6554
rect 3760 6502 3772 6554
rect 3772 6502 3786 6554
rect 3810 6502 3824 6554
rect 3824 6502 3836 6554
rect 3836 6502 3866 6554
rect 3890 6502 3900 6554
rect 3900 6502 3946 6554
rect 3650 6500 3706 6502
rect 3730 6500 3786 6502
rect 3810 6500 3866 6502
rect 3890 6500 3946 6502
rect 5006 6554 5062 6556
rect 5086 6554 5142 6556
rect 5166 6554 5222 6556
rect 5246 6554 5302 6556
rect 5006 6502 5052 6554
rect 5052 6502 5062 6554
rect 5086 6502 5116 6554
rect 5116 6502 5128 6554
rect 5128 6502 5142 6554
rect 5166 6502 5180 6554
rect 5180 6502 5192 6554
rect 5192 6502 5222 6554
rect 5246 6502 5256 6554
rect 5256 6502 5302 6554
rect 5006 6500 5062 6502
rect 5086 6500 5142 6502
rect 5166 6500 5222 6502
rect 5246 6500 5302 6502
rect 6362 6554 6418 6556
rect 6442 6554 6498 6556
rect 6522 6554 6578 6556
rect 6602 6554 6658 6556
rect 6362 6502 6408 6554
rect 6408 6502 6418 6554
rect 6442 6502 6472 6554
rect 6472 6502 6484 6554
rect 6484 6502 6498 6554
rect 6522 6502 6536 6554
rect 6536 6502 6548 6554
rect 6548 6502 6578 6554
rect 6602 6502 6612 6554
rect 6612 6502 6658 6554
rect 6362 6500 6418 6502
rect 6442 6500 6498 6502
rect 6522 6500 6578 6502
rect 6602 6500 6658 6502
rect 6182 6180 6238 6216
rect 6182 6160 6184 6180
rect 6184 6160 6236 6180
rect 6236 6160 6238 6180
rect 1634 6010 1690 6012
rect 1714 6010 1770 6012
rect 1794 6010 1850 6012
rect 1874 6010 1930 6012
rect 1634 5958 1680 6010
rect 1680 5958 1690 6010
rect 1714 5958 1744 6010
rect 1744 5958 1756 6010
rect 1756 5958 1770 6010
rect 1794 5958 1808 6010
rect 1808 5958 1820 6010
rect 1820 5958 1850 6010
rect 1874 5958 1884 6010
rect 1884 5958 1930 6010
rect 1634 5956 1690 5958
rect 1714 5956 1770 5958
rect 1794 5956 1850 5958
rect 1874 5956 1930 5958
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 3150 6010 3206 6012
rect 3230 6010 3286 6012
rect 2990 5958 3036 6010
rect 3036 5958 3046 6010
rect 3070 5958 3100 6010
rect 3100 5958 3112 6010
rect 3112 5958 3126 6010
rect 3150 5958 3164 6010
rect 3164 5958 3176 6010
rect 3176 5958 3206 6010
rect 3230 5958 3240 6010
rect 3240 5958 3286 6010
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 3150 5956 3206 5958
rect 3230 5956 3286 5958
rect 4346 6010 4402 6012
rect 4426 6010 4482 6012
rect 4506 6010 4562 6012
rect 4586 6010 4642 6012
rect 4346 5958 4392 6010
rect 4392 5958 4402 6010
rect 4426 5958 4456 6010
rect 4456 5958 4468 6010
rect 4468 5958 4482 6010
rect 4506 5958 4520 6010
rect 4520 5958 4532 6010
rect 4532 5958 4562 6010
rect 4586 5958 4596 6010
rect 4596 5958 4642 6010
rect 4346 5956 4402 5958
rect 4426 5956 4482 5958
rect 4506 5956 4562 5958
rect 4586 5956 4642 5958
rect 5702 6010 5758 6012
rect 5782 6010 5838 6012
rect 5862 6010 5918 6012
rect 5942 6010 5998 6012
rect 5702 5958 5748 6010
rect 5748 5958 5758 6010
rect 5782 5958 5812 6010
rect 5812 5958 5824 6010
rect 5824 5958 5838 6010
rect 5862 5958 5876 6010
rect 5876 5958 5888 6010
rect 5888 5958 5918 6010
rect 5942 5958 5952 6010
rect 5952 5958 5998 6010
rect 5702 5956 5758 5958
rect 5782 5956 5838 5958
rect 5862 5956 5918 5958
rect 5942 5956 5998 5958
rect 6734 5480 6790 5536
rect 2294 5466 2350 5468
rect 2374 5466 2430 5468
rect 2454 5466 2510 5468
rect 2534 5466 2590 5468
rect 2294 5414 2340 5466
rect 2340 5414 2350 5466
rect 2374 5414 2404 5466
rect 2404 5414 2416 5466
rect 2416 5414 2430 5466
rect 2454 5414 2468 5466
rect 2468 5414 2480 5466
rect 2480 5414 2510 5466
rect 2534 5414 2544 5466
rect 2544 5414 2590 5466
rect 2294 5412 2350 5414
rect 2374 5412 2430 5414
rect 2454 5412 2510 5414
rect 2534 5412 2590 5414
rect 3650 5466 3706 5468
rect 3730 5466 3786 5468
rect 3810 5466 3866 5468
rect 3890 5466 3946 5468
rect 3650 5414 3696 5466
rect 3696 5414 3706 5466
rect 3730 5414 3760 5466
rect 3760 5414 3772 5466
rect 3772 5414 3786 5466
rect 3810 5414 3824 5466
rect 3824 5414 3836 5466
rect 3836 5414 3866 5466
rect 3890 5414 3900 5466
rect 3900 5414 3946 5466
rect 3650 5412 3706 5414
rect 3730 5412 3786 5414
rect 3810 5412 3866 5414
rect 3890 5412 3946 5414
rect 5006 5466 5062 5468
rect 5086 5466 5142 5468
rect 5166 5466 5222 5468
rect 5246 5466 5302 5468
rect 5006 5414 5052 5466
rect 5052 5414 5062 5466
rect 5086 5414 5116 5466
rect 5116 5414 5128 5466
rect 5128 5414 5142 5466
rect 5166 5414 5180 5466
rect 5180 5414 5192 5466
rect 5192 5414 5222 5466
rect 5246 5414 5256 5466
rect 5256 5414 5302 5466
rect 5006 5412 5062 5414
rect 5086 5412 5142 5414
rect 5166 5412 5222 5414
rect 5246 5412 5302 5414
rect 6362 5466 6418 5468
rect 6442 5466 6498 5468
rect 6522 5466 6578 5468
rect 6602 5466 6658 5468
rect 6362 5414 6408 5466
rect 6408 5414 6418 5466
rect 6442 5414 6472 5466
rect 6472 5414 6484 5466
rect 6484 5414 6498 5466
rect 6522 5414 6536 5466
rect 6536 5414 6548 5466
rect 6548 5414 6578 5466
rect 6602 5414 6612 5466
rect 6612 5414 6658 5466
rect 6362 5412 6418 5414
rect 6442 5412 6498 5414
rect 6522 5412 6578 5414
rect 6602 5412 6658 5414
rect 1634 4922 1690 4924
rect 1714 4922 1770 4924
rect 1794 4922 1850 4924
rect 1874 4922 1930 4924
rect 1634 4870 1680 4922
rect 1680 4870 1690 4922
rect 1714 4870 1744 4922
rect 1744 4870 1756 4922
rect 1756 4870 1770 4922
rect 1794 4870 1808 4922
rect 1808 4870 1820 4922
rect 1820 4870 1850 4922
rect 1874 4870 1884 4922
rect 1884 4870 1930 4922
rect 1634 4868 1690 4870
rect 1714 4868 1770 4870
rect 1794 4868 1850 4870
rect 1874 4868 1930 4870
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 3150 4922 3206 4924
rect 3230 4922 3286 4924
rect 2990 4870 3036 4922
rect 3036 4870 3046 4922
rect 3070 4870 3100 4922
rect 3100 4870 3112 4922
rect 3112 4870 3126 4922
rect 3150 4870 3164 4922
rect 3164 4870 3176 4922
rect 3176 4870 3206 4922
rect 3230 4870 3240 4922
rect 3240 4870 3286 4922
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 3150 4868 3206 4870
rect 3230 4868 3286 4870
rect 4346 4922 4402 4924
rect 4426 4922 4482 4924
rect 4506 4922 4562 4924
rect 4586 4922 4642 4924
rect 4346 4870 4392 4922
rect 4392 4870 4402 4922
rect 4426 4870 4456 4922
rect 4456 4870 4468 4922
rect 4468 4870 4482 4922
rect 4506 4870 4520 4922
rect 4520 4870 4532 4922
rect 4532 4870 4562 4922
rect 4586 4870 4596 4922
rect 4596 4870 4642 4922
rect 4346 4868 4402 4870
rect 4426 4868 4482 4870
rect 4506 4868 4562 4870
rect 4586 4868 4642 4870
rect 5702 4922 5758 4924
rect 5782 4922 5838 4924
rect 5862 4922 5918 4924
rect 5942 4922 5998 4924
rect 5702 4870 5748 4922
rect 5748 4870 5758 4922
rect 5782 4870 5812 4922
rect 5812 4870 5824 4922
rect 5824 4870 5838 4922
rect 5862 4870 5876 4922
rect 5876 4870 5888 4922
rect 5888 4870 5918 4922
rect 5942 4870 5952 4922
rect 5952 4870 5998 4922
rect 5702 4868 5758 4870
rect 5782 4868 5838 4870
rect 5862 4868 5918 4870
rect 5942 4868 5998 4870
rect 6182 4800 6238 4856
rect 2294 4378 2350 4380
rect 2374 4378 2430 4380
rect 2454 4378 2510 4380
rect 2534 4378 2590 4380
rect 2294 4326 2340 4378
rect 2340 4326 2350 4378
rect 2374 4326 2404 4378
rect 2404 4326 2416 4378
rect 2416 4326 2430 4378
rect 2454 4326 2468 4378
rect 2468 4326 2480 4378
rect 2480 4326 2510 4378
rect 2534 4326 2544 4378
rect 2544 4326 2590 4378
rect 2294 4324 2350 4326
rect 2374 4324 2430 4326
rect 2454 4324 2510 4326
rect 2534 4324 2590 4326
rect 3650 4378 3706 4380
rect 3730 4378 3786 4380
rect 3810 4378 3866 4380
rect 3890 4378 3946 4380
rect 3650 4326 3696 4378
rect 3696 4326 3706 4378
rect 3730 4326 3760 4378
rect 3760 4326 3772 4378
rect 3772 4326 3786 4378
rect 3810 4326 3824 4378
rect 3824 4326 3836 4378
rect 3836 4326 3866 4378
rect 3890 4326 3900 4378
rect 3900 4326 3946 4378
rect 3650 4324 3706 4326
rect 3730 4324 3786 4326
rect 3810 4324 3866 4326
rect 3890 4324 3946 4326
rect 5006 4378 5062 4380
rect 5086 4378 5142 4380
rect 5166 4378 5222 4380
rect 5246 4378 5302 4380
rect 5006 4326 5052 4378
rect 5052 4326 5062 4378
rect 5086 4326 5116 4378
rect 5116 4326 5128 4378
rect 5128 4326 5142 4378
rect 5166 4326 5180 4378
rect 5180 4326 5192 4378
rect 5192 4326 5222 4378
rect 5246 4326 5256 4378
rect 5256 4326 5302 4378
rect 5006 4324 5062 4326
rect 5086 4324 5142 4326
rect 5166 4324 5222 4326
rect 5246 4324 5302 4326
rect 6362 4378 6418 4380
rect 6442 4378 6498 4380
rect 6522 4378 6578 4380
rect 6602 4378 6658 4380
rect 6362 4326 6408 4378
rect 6408 4326 6418 4378
rect 6442 4326 6472 4378
rect 6472 4326 6484 4378
rect 6484 4326 6498 4378
rect 6522 4326 6536 4378
rect 6536 4326 6548 4378
rect 6548 4326 6578 4378
rect 6602 4326 6612 4378
rect 6612 4326 6658 4378
rect 6362 4324 6418 4326
rect 6442 4324 6498 4326
rect 6522 4324 6578 4326
rect 6602 4324 6658 4326
rect 6182 4120 6238 4176
rect 1634 3834 1690 3836
rect 1714 3834 1770 3836
rect 1794 3834 1850 3836
rect 1874 3834 1930 3836
rect 1634 3782 1680 3834
rect 1680 3782 1690 3834
rect 1714 3782 1744 3834
rect 1744 3782 1756 3834
rect 1756 3782 1770 3834
rect 1794 3782 1808 3834
rect 1808 3782 1820 3834
rect 1820 3782 1850 3834
rect 1874 3782 1884 3834
rect 1884 3782 1930 3834
rect 1634 3780 1690 3782
rect 1714 3780 1770 3782
rect 1794 3780 1850 3782
rect 1874 3780 1930 3782
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 3150 3834 3206 3836
rect 3230 3834 3286 3836
rect 2990 3782 3036 3834
rect 3036 3782 3046 3834
rect 3070 3782 3100 3834
rect 3100 3782 3112 3834
rect 3112 3782 3126 3834
rect 3150 3782 3164 3834
rect 3164 3782 3176 3834
rect 3176 3782 3206 3834
rect 3230 3782 3240 3834
rect 3240 3782 3286 3834
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 3150 3780 3206 3782
rect 3230 3780 3286 3782
rect 4346 3834 4402 3836
rect 4426 3834 4482 3836
rect 4506 3834 4562 3836
rect 4586 3834 4642 3836
rect 4346 3782 4392 3834
rect 4392 3782 4402 3834
rect 4426 3782 4456 3834
rect 4456 3782 4468 3834
rect 4468 3782 4482 3834
rect 4506 3782 4520 3834
rect 4520 3782 4532 3834
rect 4532 3782 4562 3834
rect 4586 3782 4596 3834
rect 4596 3782 4642 3834
rect 4346 3780 4402 3782
rect 4426 3780 4482 3782
rect 4506 3780 4562 3782
rect 4586 3780 4642 3782
rect 5702 3834 5758 3836
rect 5782 3834 5838 3836
rect 5862 3834 5918 3836
rect 5942 3834 5998 3836
rect 5702 3782 5748 3834
rect 5748 3782 5758 3834
rect 5782 3782 5812 3834
rect 5812 3782 5824 3834
rect 5824 3782 5838 3834
rect 5862 3782 5876 3834
rect 5876 3782 5888 3834
rect 5888 3782 5918 3834
rect 5942 3782 5952 3834
rect 5952 3782 5998 3834
rect 5702 3780 5758 3782
rect 5782 3780 5838 3782
rect 5862 3780 5918 3782
rect 5942 3780 5998 3782
rect 2294 3290 2350 3292
rect 2374 3290 2430 3292
rect 2454 3290 2510 3292
rect 2534 3290 2590 3292
rect 2294 3238 2340 3290
rect 2340 3238 2350 3290
rect 2374 3238 2404 3290
rect 2404 3238 2416 3290
rect 2416 3238 2430 3290
rect 2454 3238 2468 3290
rect 2468 3238 2480 3290
rect 2480 3238 2510 3290
rect 2534 3238 2544 3290
rect 2544 3238 2590 3290
rect 2294 3236 2350 3238
rect 2374 3236 2430 3238
rect 2454 3236 2510 3238
rect 2534 3236 2590 3238
rect 3650 3290 3706 3292
rect 3730 3290 3786 3292
rect 3810 3290 3866 3292
rect 3890 3290 3946 3292
rect 3650 3238 3696 3290
rect 3696 3238 3706 3290
rect 3730 3238 3760 3290
rect 3760 3238 3772 3290
rect 3772 3238 3786 3290
rect 3810 3238 3824 3290
rect 3824 3238 3836 3290
rect 3836 3238 3866 3290
rect 3890 3238 3900 3290
rect 3900 3238 3946 3290
rect 3650 3236 3706 3238
rect 3730 3236 3786 3238
rect 3810 3236 3866 3238
rect 3890 3236 3946 3238
rect 5006 3290 5062 3292
rect 5086 3290 5142 3292
rect 5166 3290 5222 3292
rect 5246 3290 5302 3292
rect 5006 3238 5052 3290
rect 5052 3238 5062 3290
rect 5086 3238 5116 3290
rect 5116 3238 5128 3290
rect 5128 3238 5142 3290
rect 5166 3238 5180 3290
rect 5180 3238 5192 3290
rect 5192 3238 5222 3290
rect 5246 3238 5256 3290
rect 5256 3238 5302 3290
rect 5006 3236 5062 3238
rect 5086 3236 5142 3238
rect 5166 3236 5222 3238
rect 5246 3236 5302 3238
rect 6362 3290 6418 3292
rect 6442 3290 6498 3292
rect 6522 3290 6578 3292
rect 6602 3290 6658 3292
rect 6362 3238 6408 3290
rect 6408 3238 6418 3290
rect 6442 3238 6472 3290
rect 6472 3238 6484 3290
rect 6484 3238 6498 3290
rect 6522 3238 6536 3290
rect 6536 3238 6548 3290
rect 6548 3238 6578 3290
rect 6602 3238 6612 3290
rect 6612 3238 6658 3290
rect 6362 3236 6418 3238
rect 6442 3236 6498 3238
rect 6522 3236 6578 3238
rect 6602 3236 6658 3238
rect 1634 2746 1690 2748
rect 1714 2746 1770 2748
rect 1794 2746 1850 2748
rect 1874 2746 1930 2748
rect 1634 2694 1680 2746
rect 1680 2694 1690 2746
rect 1714 2694 1744 2746
rect 1744 2694 1756 2746
rect 1756 2694 1770 2746
rect 1794 2694 1808 2746
rect 1808 2694 1820 2746
rect 1820 2694 1850 2746
rect 1874 2694 1884 2746
rect 1884 2694 1930 2746
rect 1634 2692 1690 2694
rect 1714 2692 1770 2694
rect 1794 2692 1850 2694
rect 1874 2692 1930 2694
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 3150 2746 3206 2748
rect 3230 2746 3286 2748
rect 2990 2694 3036 2746
rect 3036 2694 3046 2746
rect 3070 2694 3100 2746
rect 3100 2694 3112 2746
rect 3112 2694 3126 2746
rect 3150 2694 3164 2746
rect 3164 2694 3176 2746
rect 3176 2694 3206 2746
rect 3230 2694 3240 2746
rect 3240 2694 3286 2746
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 3150 2692 3206 2694
rect 3230 2692 3286 2694
rect 4346 2746 4402 2748
rect 4426 2746 4482 2748
rect 4506 2746 4562 2748
rect 4586 2746 4642 2748
rect 4346 2694 4392 2746
rect 4392 2694 4402 2746
rect 4426 2694 4456 2746
rect 4456 2694 4468 2746
rect 4468 2694 4482 2746
rect 4506 2694 4520 2746
rect 4520 2694 4532 2746
rect 4532 2694 4562 2746
rect 4586 2694 4596 2746
rect 4596 2694 4642 2746
rect 4346 2692 4402 2694
rect 4426 2692 4482 2694
rect 4506 2692 4562 2694
rect 4586 2692 4642 2694
rect 5702 2746 5758 2748
rect 5782 2746 5838 2748
rect 5862 2746 5918 2748
rect 5942 2746 5998 2748
rect 5702 2694 5748 2746
rect 5748 2694 5758 2746
rect 5782 2694 5812 2746
rect 5812 2694 5824 2746
rect 5824 2694 5838 2746
rect 5862 2694 5876 2746
rect 5876 2694 5888 2746
rect 5888 2694 5918 2746
rect 5942 2694 5952 2746
rect 5952 2694 5998 2746
rect 5702 2692 5758 2694
rect 5782 2692 5838 2694
rect 5862 2692 5918 2694
rect 5942 2692 5998 2694
rect 2294 2202 2350 2204
rect 2374 2202 2430 2204
rect 2454 2202 2510 2204
rect 2534 2202 2590 2204
rect 2294 2150 2340 2202
rect 2340 2150 2350 2202
rect 2374 2150 2404 2202
rect 2404 2150 2416 2202
rect 2416 2150 2430 2202
rect 2454 2150 2468 2202
rect 2468 2150 2480 2202
rect 2480 2150 2510 2202
rect 2534 2150 2544 2202
rect 2544 2150 2590 2202
rect 2294 2148 2350 2150
rect 2374 2148 2430 2150
rect 2454 2148 2510 2150
rect 2534 2148 2590 2150
rect 3650 2202 3706 2204
rect 3730 2202 3786 2204
rect 3810 2202 3866 2204
rect 3890 2202 3946 2204
rect 3650 2150 3696 2202
rect 3696 2150 3706 2202
rect 3730 2150 3760 2202
rect 3760 2150 3772 2202
rect 3772 2150 3786 2202
rect 3810 2150 3824 2202
rect 3824 2150 3836 2202
rect 3836 2150 3866 2202
rect 3890 2150 3900 2202
rect 3900 2150 3946 2202
rect 3650 2148 3706 2150
rect 3730 2148 3786 2150
rect 3810 2148 3866 2150
rect 3890 2148 3946 2150
rect 5006 2202 5062 2204
rect 5086 2202 5142 2204
rect 5166 2202 5222 2204
rect 5246 2202 5302 2204
rect 5006 2150 5052 2202
rect 5052 2150 5062 2202
rect 5086 2150 5116 2202
rect 5116 2150 5128 2202
rect 5128 2150 5142 2202
rect 5166 2150 5180 2202
rect 5180 2150 5192 2202
rect 5192 2150 5222 2202
rect 5246 2150 5256 2202
rect 5256 2150 5302 2202
rect 5006 2148 5062 2150
rect 5086 2148 5142 2150
rect 5166 2148 5222 2150
rect 5246 2148 5302 2150
rect 6362 2202 6418 2204
rect 6442 2202 6498 2204
rect 6522 2202 6578 2204
rect 6602 2202 6658 2204
rect 6362 2150 6408 2202
rect 6408 2150 6418 2202
rect 6442 2150 6472 2202
rect 6472 2150 6484 2202
rect 6484 2150 6498 2202
rect 6522 2150 6536 2202
rect 6536 2150 6548 2202
rect 6548 2150 6578 2202
rect 6602 2150 6612 2202
rect 6612 2150 6658 2202
rect 6362 2148 6418 2150
rect 6442 2148 6498 2150
rect 6522 2148 6578 2150
rect 6602 2148 6658 2150
<< metal3 >>
rect 2284 7648 2600 7649
rect 2284 7584 2290 7648
rect 2354 7584 2370 7648
rect 2434 7584 2450 7648
rect 2514 7584 2530 7648
rect 2594 7584 2600 7648
rect 2284 7583 2600 7584
rect 3640 7648 3956 7649
rect 3640 7584 3646 7648
rect 3710 7584 3726 7648
rect 3790 7584 3806 7648
rect 3870 7584 3886 7648
rect 3950 7584 3956 7648
rect 3640 7583 3956 7584
rect 4996 7648 5312 7649
rect 4996 7584 5002 7648
rect 5066 7584 5082 7648
rect 5146 7584 5162 7648
rect 5226 7584 5242 7648
rect 5306 7584 5312 7648
rect 4996 7583 5312 7584
rect 6352 7648 6668 7649
rect 6352 7584 6358 7648
rect 6422 7584 6438 7648
rect 6502 7584 6518 7648
rect 6582 7584 6598 7648
rect 6662 7584 6668 7648
rect 6352 7583 6668 7584
rect 1624 7104 1940 7105
rect 1624 7040 1630 7104
rect 1694 7040 1710 7104
rect 1774 7040 1790 7104
rect 1854 7040 1870 7104
rect 1934 7040 1940 7104
rect 1624 7039 1940 7040
rect 2980 7104 3296 7105
rect 2980 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3146 7104
rect 3210 7040 3226 7104
rect 3290 7040 3296 7104
rect 2980 7039 3296 7040
rect 4336 7104 4652 7105
rect 4336 7040 4342 7104
rect 4406 7040 4422 7104
rect 4486 7040 4502 7104
rect 4566 7040 4582 7104
rect 4646 7040 4652 7104
rect 4336 7039 4652 7040
rect 5692 7104 6008 7105
rect 5692 7040 5698 7104
rect 5762 7040 5778 7104
rect 5842 7040 5858 7104
rect 5922 7040 5938 7104
rect 6002 7040 6008 7104
rect 5692 7039 6008 7040
rect 2284 6560 2600 6561
rect 2284 6496 2290 6560
rect 2354 6496 2370 6560
rect 2434 6496 2450 6560
rect 2514 6496 2530 6560
rect 2594 6496 2600 6560
rect 2284 6495 2600 6496
rect 3640 6560 3956 6561
rect 3640 6496 3646 6560
rect 3710 6496 3726 6560
rect 3790 6496 3806 6560
rect 3870 6496 3886 6560
rect 3950 6496 3956 6560
rect 3640 6495 3956 6496
rect 4996 6560 5312 6561
rect 4996 6496 5002 6560
rect 5066 6496 5082 6560
rect 5146 6496 5162 6560
rect 5226 6496 5242 6560
rect 5306 6496 5312 6560
rect 4996 6495 5312 6496
rect 6352 6560 6668 6561
rect 6352 6496 6358 6560
rect 6422 6496 6438 6560
rect 6502 6496 6518 6560
rect 6582 6496 6598 6560
rect 6662 6496 6668 6560
rect 6352 6495 6668 6496
rect 6177 6218 6243 6221
rect 6888 6218 7688 6248
rect 6177 6216 7688 6218
rect 6177 6160 6182 6216
rect 6238 6160 7688 6216
rect 6177 6158 7688 6160
rect 6177 6155 6243 6158
rect 6888 6128 7688 6158
rect 1624 6016 1940 6017
rect 1624 5952 1630 6016
rect 1694 5952 1710 6016
rect 1774 5952 1790 6016
rect 1854 5952 1870 6016
rect 1934 5952 1940 6016
rect 1624 5951 1940 5952
rect 2980 6016 3296 6017
rect 2980 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3146 6016
rect 3210 5952 3226 6016
rect 3290 5952 3296 6016
rect 2980 5951 3296 5952
rect 4336 6016 4652 6017
rect 4336 5952 4342 6016
rect 4406 5952 4422 6016
rect 4486 5952 4502 6016
rect 4566 5952 4582 6016
rect 4646 5952 4652 6016
rect 4336 5951 4652 5952
rect 5692 6016 6008 6017
rect 5692 5952 5698 6016
rect 5762 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5938 6016
rect 6002 5952 6008 6016
rect 5692 5951 6008 5952
rect 6729 5538 6795 5541
rect 6888 5538 7688 5568
rect 6729 5536 7688 5538
rect 6729 5480 6734 5536
rect 6790 5480 7688 5536
rect 6729 5478 7688 5480
rect 6729 5475 6795 5478
rect 2284 5472 2600 5473
rect 2284 5408 2290 5472
rect 2354 5408 2370 5472
rect 2434 5408 2450 5472
rect 2514 5408 2530 5472
rect 2594 5408 2600 5472
rect 2284 5407 2600 5408
rect 3640 5472 3956 5473
rect 3640 5408 3646 5472
rect 3710 5408 3726 5472
rect 3790 5408 3806 5472
rect 3870 5408 3886 5472
rect 3950 5408 3956 5472
rect 3640 5407 3956 5408
rect 4996 5472 5312 5473
rect 4996 5408 5002 5472
rect 5066 5408 5082 5472
rect 5146 5408 5162 5472
rect 5226 5408 5242 5472
rect 5306 5408 5312 5472
rect 4996 5407 5312 5408
rect 6352 5472 6668 5473
rect 6352 5408 6358 5472
rect 6422 5408 6438 5472
rect 6502 5408 6518 5472
rect 6582 5408 6598 5472
rect 6662 5408 6668 5472
rect 6888 5448 7688 5478
rect 6352 5407 6668 5408
rect 1624 4928 1940 4929
rect 1624 4864 1630 4928
rect 1694 4864 1710 4928
rect 1774 4864 1790 4928
rect 1854 4864 1870 4928
rect 1934 4864 1940 4928
rect 1624 4863 1940 4864
rect 2980 4928 3296 4929
rect 2980 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3146 4928
rect 3210 4864 3226 4928
rect 3290 4864 3296 4928
rect 2980 4863 3296 4864
rect 4336 4928 4652 4929
rect 4336 4864 4342 4928
rect 4406 4864 4422 4928
rect 4486 4864 4502 4928
rect 4566 4864 4582 4928
rect 4646 4864 4652 4928
rect 4336 4863 4652 4864
rect 5692 4928 6008 4929
rect 5692 4864 5698 4928
rect 5762 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5938 4928
rect 6002 4864 6008 4928
rect 5692 4863 6008 4864
rect 6177 4858 6243 4861
rect 6888 4858 7688 4888
rect 6177 4856 7688 4858
rect 6177 4800 6182 4856
rect 6238 4800 7688 4856
rect 6177 4798 7688 4800
rect 6177 4795 6243 4798
rect 6888 4768 7688 4798
rect 2284 4384 2600 4385
rect 2284 4320 2290 4384
rect 2354 4320 2370 4384
rect 2434 4320 2450 4384
rect 2514 4320 2530 4384
rect 2594 4320 2600 4384
rect 2284 4319 2600 4320
rect 3640 4384 3956 4385
rect 3640 4320 3646 4384
rect 3710 4320 3726 4384
rect 3790 4320 3806 4384
rect 3870 4320 3886 4384
rect 3950 4320 3956 4384
rect 3640 4319 3956 4320
rect 4996 4384 5312 4385
rect 4996 4320 5002 4384
rect 5066 4320 5082 4384
rect 5146 4320 5162 4384
rect 5226 4320 5242 4384
rect 5306 4320 5312 4384
rect 4996 4319 5312 4320
rect 6352 4384 6668 4385
rect 6352 4320 6358 4384
rect 6422 4320 6438 4384
rect 6502 4320 6518 4384
rect 6582 4320 6598 4384
rect 6662 4320 6668 4384
rect 6352 4319 6668 4320
rect 6177 4178 6243 4181
rect 6888 4178 7688 4208
rect 6177 4176 7688 4178
rect 6177 4120 6182 4176
rect 6238 4120 7688 4176
rect 6177 4118 7688 4120
rect 6177 4115 6243 4118
rect 6888 4088 7688 4118
rect 1624 3840 1940 3841
rect 1624 3776 1630 3840
rect 1694 3776 1710 3840
rect 1774 3776 1790 3840
rect 1854 3776 1870 3840
rect 1934 3776 1940 3840
rect 1624 3775 1940 3776
rect 2980 3840 3296 3841
rect 2980 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3146 3840
rect 3210 3776 3226 3840
rect 3290 3776 3296 3840
rect 2980 3775 3296 3776
rect 4336 3840 4652 3841
rect 4336 3776 4342 3840
rect 4406 3776 4422 3840
rect 4486 3776 4502 3840
rect 4566 3776 4582 3840
rect 4646 3776 4652 3840
rect 4336 3775 4652 3776
rect 5692 3840 6008 3841
rect 5692 3776 5698 3840
rect 5762 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5938 3840
rect 6002 3776 6008 3840
rect 5692 3775 6008 3776
rect 2284 3296 2600 3297
rect 2284 3232 2290 3296
rect 2354 3232 2370 3296
rect 2434 3232 2450 3296
rect 2514 3232 2530 3296
rect 2594 3232 2600 3296
rect 2284 3231 2600 3232
rect 3640 3296 3956 3297
rect 3640 3232 3646 3296
rect 3710 3232 3726 3296
rect 3790 3232 3806 3296
rect 3870 3232 3886 3296
rect 3950 3232 3956 3296
rect 3640 3231 3956 3232
rect 4996 3296 5312 3297
rect 4996 3232 5002 3296
rect 5066 3232 5082 3296
rect 5146 3232 5162 3296
rect 5226 3232 5242 3296
rect 5306 3232 5312 3296
rect 4996 3231 5312 3232
rect 6352 3296 6668 3297
rect 6352 3232 6358 3296
rect 6422 3232 6438 3296
rect 6502 3232 6518 3296
rect 6582 3232 6598 3296
rect 6662 3232 6668 3296
rect 6352 3231 6668 3232
rect 1624 2752 1940 2753
rect 1624 2688 1630 2752
rect 1694 2688 1710 2752
rect 1774 2688 1790 2752
rect 1854 2688 1870 2752
rect 1934 2688 1940 2752
rect 1624 2687 1940 2688
rect 2980 2752 3296 2753
rect 2980 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3146 2752
rect 3210 2688 3226 2752
rect 3290 2688 3296 2752
rect 2980 2687 3296 2688
rect 4336 2752 4652 2753
rect 4336 2688 4342 2752
rect 4406 2688 4422 2752
rect 4486 2688 4502 2752
rect 4566 2688 4582 2752
rect 4646 2688 4652 2752
rect 4336 2687 4652 2688
rect 5692 2752 6008 2753
rect 5692 2688 5698 2752
rect 5762 2688 5778 2752
rect 5842 2688 5858 2752
rect 5922 2688 5938 2752
rect 6002 2688 6008 2752
rect 5692 2687 6008 2688
rect 2284 2208 2600 2209
rect 2284 2144 2290 2208
rect 2354 2144 2370 2208
rect 2434 2144 2450 2208
rect 2514 2144 2530 2208
rect 2594 2144 2600 2208
rect 2284 2143 2600 2144
rect 3640 2208 3956 2209
rect 3640 2144 3646 2208
rect 3710 2144 3726 2208
rect 3790 2144 3806 2208
rect 3870 2144 3886 2208
rect 3950 2144 3956 2208
rect 3640 2143 3956 2144
rect 4996 2208 5312 2209
rect 4996 2144 5002 2208
rect 5066 2144 5082 2208
rect 5146 2144 5162 2208
rect 5226 2144 5242 2208
rect 5306 2144 5312 2208
rect 4996 2143 5312 2144
rect 6352 2208 6668 2209
rect 6352 2144 6358 2208
rect 6422 2144 6438 2208
rect 6502 2144 6518 2208
rect 6582 2144 6598 2208
rect 6662 2144 6668 2208
rect 6352 2143 6668 2144
<< via3 >>
rect 2290 7644 2354 7648
rect 2290 7588 2294 7644
rect 2294 7588 2350 7644
rect 2350 7588 2354 7644
rect 2290 7584 2354 7588
rect 2370 7644 2434 7648
rect 2370 7588 2374 7644
rect 2374 7588 2430 7644
rect 2430 7588 2434 7644
rect 2370 7584 2434 7588
rect 2450 7644 2514 7648
rect 2450 7588 2454 7644
rect 2454 7588 2510 7644
rect 2510 7588 2514 7644
rect 2450 7584 2514 7588
rect 2530 7644 2594 7648
rect 2530 7588 2534 7644
rect 2534 7588 2590 7644
rect 2590 7588 2594 7644
rect 2530 7584 2594 7588
rect 3646 7644 3710 7648
rect 3646 7588 3650 7644
rect 3650 7588 3706 7644
rect 3706 7588 3710 7644
rect 3646 7584 3710 7588
rect 3726 7644 3790 7648
rect 3726 7588 3730 7644
rect 3730 7588 3786 7644
rect 3786 7588 3790 7644
rect 3726 7584 3790 7588
rect 3806 7644 3870 7648
rect 3806 7588 3810 7644
rect 3810 7588 3866 7644
rect 3866 7588 3870 7644
rect 3806 7584 3870 7588
rect 3886 7644 3950 7648
rect 3886 7588 3890 7644
rect 3890 7588 3946 7644
rect 3946 7588 3950 7644
rect 3886 7584 3950 7588
rect 5002 7644 5066 7648
rect 5002 7588 5006 7644
rect 5006 7588 5062 7644
rect 5062 7588 5066 7644
rect 5002 7584 5066 7588
rect 5082 7644 5146 7648
rect 5082 7588 5086 7644
rect 5086 7588 5142 7644
rect 5142 7588 5146 7644
rect 5082 7584 5146 7588
rect 5162 7644 5226 7648
rect 5162 7588 5166 7644
rect 5166 7588 5222 7644
rect 5222 7588 5226 7644
rect 5162 7584 5226 7588
rect 5242 7644 5306 7648
rect 5242 7588 5246 7644
rect 5246 7588 5302 7644
rect 5302 7588 5306 7644
rect 5242 7584 5306 7588
rect 6358 7644 6422 7648
rect 6358 7588 6362 7644
rect 6362 7588 6418 7644
rect 6418 7588 6422 7644
rect 6358 7584 6422 7588
rect 6438 7644 6502 7648
rect 6438 7588 6442 7644
rect 6442 7588 6498 7644
rect 6498 7588 6502 7644
rect 6438 7584 6502 7588
rect 6518 7644 6582 7648
rect 6518 7588 6522 7644
rect 6522 7588 6578 7644
rect 6578 7588 6582 7644
rect 6518 7584 6582 7588
rect 6598 7644 6662 7648
rect 6598 7588 6602 7644
rect 6602 7588 6658 7644
rect 6658 7588 6662 7644
rect 6598 7584 6662 7588
rect 1630 7100 1694 7104
rect 1630 7044 1634 7100
rect 1634 7044 1690 7100
rect 1690 7044 1694 7100
rect 1630 7040 1694 7044
rect 1710 7100 1774 7104
rect 1710 7044 1714 7100
rect 1714 7044 1770 7100
rect 1770 7044 1774 7100
rect 1710 7040 1774 7044
rect 1790 7100 1854 7104
rect 1790 7044 1794 7100
rect 1794 7044 1850 7100
rect 1850 7044 1854 7100
rect 1790 7040 1854 7044
rect 1870 7100 1934 7104
rect 1870 7044 1874 7100
rect 1874 7044 1930 7100
rect 1930 7044 1934 7100
rect 1870 7040 1934 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 3146 7100 3210 7104
rect 3146 7044 3150 7100
rect 3150 7044 3206 7100
rect 3206 7044 3210 7100
rect 3146 7040 3210 7044
rect 3226 7100 3290 7104
rect 3226 7044 3230 7100
rect 3230 7044 3286 7100
rect 3286 7044 3290 7100
rect 3226 7040 3290 7044
rect 4342 7100 4406 7104
rect 4342 7044 4346 7100
rect 4346 7044 4402 7100
rect 4402 7044 4406 7100
rect 4342 7040 4406 7044
rect 4422 7100 4486 7104
rect 4422 7044 4426 7100
rect 4426 7044 4482 7100
rect 4482 7044 4486 7100
rect 4422 7040 4486 7044
rect 4502 7100 4566 7104
rect 4502 7044 4506 7100
rect 4506 7044 4562 7100
rect 4562 7044 4566 7100
rect 4502 7040 4566 7044
rect 4582 7100 4646 7104
rect 4582 7044 4586 7100
rect 4586 7044 4642 7100
rect 4642 7044 4646 7100
rect 4582 7040 4646 7044
rect 5698 7100 5762 7104
rect 5698 7044 5702 7100
rect 5702 7044 5758 7100
rect 5758 7044 5762 7100
rect 5698 7040 5762 7044
rect 5778 7100 5842 7104
rect 5778 7044 5782 7100
rect 5782 7044 5838 7100
rect 5838 7044 5842 7100
rect 5778 7040 5842 7044
rect 5858 7100 5922 7104
rect 5858 7044 5862 7100
rect 5862 7044 5918 7100
rect 5918 7044 5922 7100
rect 5858 7040 5922 7044
rect 5938 7100 6002 7104
rect 5938 7044 5942 7100
rect 5942 7044 5998 7100
rect 5998 7044 6002 7100
rect 5938 7040 6002 7044
rect 2290 6556 2354 6560
rect 2290 6500 2294 6556
rect 2294 6500 2350 6556
rect 2350 6500 2354 6556
rect 2290 6496 2354 6500
rect 2370 6556 2434 6560
rect 2370 6500 2374 6556
rect 2374 6500 2430 6556
rect 2430 6500 2434 6556
rect 2370 6496 2434 6500
rect 2450 6556 2514 6560
rect 2450 6500 2454 6556
rect 2454 6500 2510 6556
rect 2510 6500 2514 6556
rect 2450 6496 2514 6500
rect 2530 6556 2594 6560
rect 2530 6500 2534 6556
rect 2534 6500 2590 6556
rect 2590 6500 2594 6556
rect 2530 6496 2594 6500
rect 3646 6556 3710 6560
rect 3646 6500 3650 6556
rect 3650 6500 3706 6556
rect 3706 6500 3710 6556
rect 3646 6496 3710 6500
rect 3726 6556 3790 6560
rect 3726 6500 3730 6556
rect 3730 6500 3786 6556
rect 3786 6500 3790 6556
rect 3726 6496 3790 6500
rect 3806 6556 3870 6560
rect 3806 6500 3810 6556
rect 3810 6500 3866 6556
rect 3866 6500 3870 6556
rect 3806 6496 3870 6500
rect 3886 6556 3950 6560
rect 3886 6500 3890 6556
rect 3890 6500 3946 6556
rect 3946 6500 3950 6556
rect 3886 6496 3950 6500
rect 5002 6556 5066 6560
rect 5002 6500 5006 6556
rect 5006 6500 5062 6556
rect 5062 6500 5066 6556
rect 5002 6496 5066 6500
rect 5082 6556 5146 6560
rect 5082 6500 5086 6556
rect 5086 6500 5142 6556
rect 5142 6500 5146 6556
rect 5082 6496 5146 6500
rect 5162 6556 5226 6560
rect 5162 6500 5166 6556
rect 5166 6500 5222 6556
rect 5222 6500 5226 6556
rect 5162 6496 5226 6500
rect 5242 6556 5306 6560
rect 5242 6500 5246 6556
rect 5246 6500 5302 6556
rect 5302 6500 5306 6556
rect 5242 6496 5306 6500
rect 6358 6556 6422 6560
rect 6358 6500 6362 6556
rect 6362 6500 6418 6556
rect 6418 6500 6422 6556
rect 6358 6496 6422 6500
rect 6438 6556 6502 6560
rect 6438 6500 6442 6556
rect 6442 6500 6498 6556
rect 6498 6500 6502 6556
rect 6438 6496 6502 6500
rect 6518 6556 6582 6560
rect 6518 6500 6522 6556
rect 6522 6500 6578 6556
rect 6578 6500 6582 6556
rect 6518 6496 6582 6500
rect 6598 6556 6662 6560
rect 6598 6500 6602 6556
rect 6602 6500 6658 6556
rect 6658 6500 6662 6556
rect 6598 6496 6662 6500
rect 1630 6012 1694 6016
rect 1630 5956 1634 6012
rect 1634 5956 1690 6012
rect 1690 5956 1694 6012
rect 1630 5952 1694 5956
rect 1710 6012 1774 6016
rect 1710 5956 1714 6012
rect 1714 5956 1770 6012
rect 1770 5956 1774 6012
rect 1710 5952 1774 5956
rect 1790 6012 1854 6016
rect 1790 5956 1794 6012
rect 1794 5956 1850 6012
rect 1850 5956 1854 6012
rect 1790 5952 1854 5956
rect 1870 6012 1934 6016
rect 1870 5956 1874 6012
rect 1874 5956 1930 6012
rect 1930 5956 1934 6012
rect 1870 5952 1934 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 3146 6012 3210 6016
rect 3146 5956 3150 6012
rect 3150 5956 3206 6012
rect 3206 5956 3210 6012
rect 3146 5952 3210 5956
rect 3226 6012 3290 6016
rect 3226 5956 3230 6012
rect 3230 5956 3286 6012
rect 3286 5956 3290 6012
rect 3226 5952 3290 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 4422 6012 4486 6016
rect 4422 5956 4426 6012
rect 4426 5956 4482 6012
rect 4482 5956 4486 6012
rect 4422 5952 4486 5956
rect 4502 6012 4566 6016
rect 4502 5956 4506 6012
rect 4506 5956 4562 6012
rect 4562 5956 4566 6012
rect 4502 5952 4566 5956
rect 4582 6012 4646 6016
rect 4582 5956 4586 6012
rect 4586 5956 4642 6012
rect 4642 5956 4646 6012
rect 4582 5952 4646 5956
rect 5698 6012 5762 6016
rect 5698 5956 5702 6012
rect 5702 5956 5758 6012
rect 5758 5956 5762 6012
rect 5698 5952 5762 5956
rect 5778 6012 5842 6016
rect 5778 5956 5782 6012
rect 5782 5956 5838 6012
rect 5838 5956 5842 6012
rect 5778 5952 5842 5956
rect 5858 6012 5922 6016
rect 5858 5956 5862 6012
rect 5862 5956 5918 6012
rect 5918 5956 5922 6012
rect 5858 5952 5922 5956
rect 5938 6012 6002 6016
rect 5938 5956 5942 6012
rect 5942 5956 5998 6012
rect 5998 5956 6002 6012
rect 5938 5952 6002 5956
rect 2290 5468 2354 5472
rect 2290 5412 2294 5468
rect 2294 5412 2350 5468
rect 2350 5412 2354 5468
rect 2290 5408 2354 5412
rect 2370 5468 2434 5472
rect 2370 5412 2374 5468
rect 2374 5412 2430 5468
rect 2430 5412 2434 5468
rect 2370 5408 2434 5412
rect 2450 5468 2514 5472
rect 2450 5412 2454 5468
rect 2454 5412 2510 5468
rect 2510 5412 2514 5468
rect 2450 5408 2514 5412
rect 2530 5468 2594 5472
rect 2530 5412 2534 5468
rect 2534 5412 2590 5468
rect 2590 5412 2594 5468
rect 2530 5408 2594 5412
rect 3646 5468 3710 5472
rect 3646 5412 3650 5468
rect 3650 5412 3706 5468
rect 3706 5412 3710 5468
rect 3646 5408 3710 5412
rect 3726 5468 3790 5472
rect 3726 5412 3730 5468
rect 3730 5412 3786 5468
rect 3786 5412 3790 5468
rect 3726 5408 3790 5412
rect 3806 5468 3870 5472
rect 3806 5412 3810 5468
rect 3810 5412 3866 5468
rect 3866 5412 3870 5468
rect 3806 5408 3870 5412
rect 3886 5468 3950 5472
rect 3886 5412 3890 5468
rect 3890 5412 3946 5468
rect 3946 5412 3950 5468
rect 3886 5408 3950 5412
rect 5002 5468 5066 5472
rect 5002 5412 5006 5468
rect 5006 5412 5062 5468
rect 5062 5412 5066 5468
rect 5002 5408 5066 5412
rect 5082 5468 5146 5472
rect 5082 5412 5086 5468
rect 5086 5412 5142 5468
rect 5142 5412 5146 5468
rect 5082 5408 5146 5412
rect 5162 5468 5226 5472
rect 5162 5412 5166 5468
rect 5166 5412 5222 5468
rect 5222 5412 5226 5468
rect 5162 5408 5226 5412
rect 5242 5468 5306 5472
rect 5242 5412 5246 5468
rect 5246 5412 5302 5468
rect 5302 5412 5306 5468
rect 5242 5408 5306 5412
rect 6358 5468 6422 5472
rect 6358 5412 6362 5468
rect 6362 5412 6418 5468
rect 6418 5412 6422 5468
rect 6358 5408 6422 5412
rect 6438 5468 6502 5472
rect 6438 5412 6442 5468
rect 6442 5412 6498 5468
rect 6498 5412 6502 5468
rect 6438 5408 6502 5412
rect 6518 5468 6582 5472
rect 6518 5412 6522 5468
rect 6522 5412 6578 5468
rect 6578 5412 6582 5468
rect 6518 5408 6582 5412
rect 6598 5468 6662 5472
rect 6598 5412 6602 5468
rect 6602 5412 6658 5468
rect 6658 5412 6662 5468
rect 6598 5408 6662 5412
rect 1630 4924 1694 4928
rect 1630 4868 1634 4924
rect 1634 4868 1690 4924
rect 1690 4868 1694 4924
rect 1630 4864 1694 4868
rect 1710 4924 1774 4928
rect 1710 4868 1714 4924
rect 1714 4868 1770 4924
rect 1770 4868 1774 4924
rect 1710 4864 1774 4868
rect 1790 4924 1854 4928
rect 1790 4868 1794 4924
rect 1794 4868 1850 4924
rect 1850 4868 1854 4924
rect 1790 4864 1854 4868
rect 1870 4924 1934 4928
rect 1870 4868 1874 4924
rect 1874 4868 1930 4924
rect 1930 4868 1934 4924
rect 1870 4864 1934 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 3146 4924 3210 4928
rect 3146 4868 3150 4924
rect 3150 4868 3206 4924
rect 3206 4868 3210 4924
rect 3146 4864 3210 4868
rect 3226 4924 3290 4928
rect 3226 4868 3230 4924
rect 3230 4868 3286 4924
rect 3286 4868 3290 4924
rect 3226 4864 3290 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 4422 4924 4486 4928
rect 4422 4868 4426 4924
rect 4426 4868 4482 4924
rect 4482 4868 4486 4924
rect 4422 4864 4486 4868
rect 4502 4924 4566 4928
rect 4502 4868 4506 4924
rect 4506 4868 4562 4924
rect 4562 4868 4566 4924
rect 4502 4864 4566 4868
rect 4582 4924 4646 4928
rect 4582 4868 4586 4924
rect 4586 4868 4642 4924
rect 4642 4868 4646 4924
rect 4582 4864 4646 4868
rect 5698 4924 5762 4928
rect 5698 4868 5702 4924
rect 5702 4868 5758 4924
rect 5758 4868 5762 4924
rect 5698 4864 5762 4868
rect 5778 4924 5842 4928
rect 5778 4868 5782 4924
rect 5782 4868 5838 4924
rect 5838 4868 5842 4924
rect 5778 4864 5842 4868
rect 5858 4924 5922 4928
rect 5858 4868 5862 4924
rect 5862 4868 5918 4924
rect 5918 4868 5922 4924
rect 5858 4864 5922 4868
rect 5938 4924 6002 4928
rect 5938 4868 5942 4924
rect 5942 4868 5998 4924
rect 5998 4868 6002 4924
rect 5938 4864 6002 4868
rect 2290 4380 2354 4384
rect 2290 4324 2294 4380
rect 2294 4324 2350 4380
rect 2350 4324 2354 4380
rect 2290 4320 2354 4324
rect 2370 4380 2434 4384
rect 2370 4324 2374 4380
rect 2374 4324 2430 4380
rect 2430 4324 2434 4380
rect 2370 4320 2434 4324
rect 2450 4380 2514 4384
rect 2450 4324 2454 4380
rect 2454 4324 2510 4380
rect 2510 4324 2514 4380
rect 2450 4320 2514 4324
rect 2530 4380 2594 4384
rect 2530 4324 2534 4380
rect 2534 4324 2590 4380
rect 2590 4324 2594 4380
rect 2530 4320 2594 4324
rect 3646 4380 3710 4384
rect 3646 4324 3650 4380
rect 3650 4324 3706 4380
rect 3706 4324 3710 4380
rect 3646 4320 3710 4324
rect 3726 4380 3790 4384
rect 3726 4324 3730 4380
rect 3730 4324 3786 4380
rect 3786 4324 3790 4380
rect 3726 4320 3790 4324
rect 3806 4380 3870 4384
rect 3806 4324 3810 4380
rect 3810 4324 3866 4380
rect 3866 4324 3870 4380
rect 3806 4320 3870 4324
rect 3886 4380 3950 4384
rect 3886 4324 3890 4380
rect 3890 4324 3946 4380
rect 3946 4324 3950 4380
rect 3886 4320 3950 4324
rect 5002 4380 5066 4384
rect 5002 4324 5006 4380
rect 5006 4324 5062 4380
rect 5062 4324 5066 4380
rect 5002 4320 5066 4324
rect 5082 4380 5146 4384
rect 5082 4324 5086 4380
rect 5086 4324 5142 4380
rect 5142 4324 5146 4380
rect 5082 4320 5146 4324
rect 5162 4380 5226 4384
rect 5162 4324 5166 4380
rect 5166 4324 5222 4380
rect 5222 4324 5226 4380
rect 5162 4320 5226 4324
rect 5242 4380 5306 4384
rect 5242 4324 5246 4380
rect 5246 4324 5302 4380
rect 5302 4324 5306 4380
rect 5242 4320 5306 4324
rect 6358 4380 6422 4384
rect 6358 4324 6362 4380
rect 6362 4324 6418 4380
rect 6418 4324 6422 4380
rect 6358 4320 6422 4324
rect 6438 4380 6502 4384
rect 6438 4324 6442 4380
rect 6442 4324 6498 4380
rect 6498 4324 6502 4380
rect 6438 4320 6502 4324
rect 6518 4380 6582 4384
rect 6518 4324 6522 4380
rect 6522 4324 6578 4380
rect 6578 4324 6582 4380
rect 6518 4320 6582 4324
rect 6598 4380 6662 4384
rect 6598 4324 6602 4380
rect 6602 4324 6658 4380
rect 6658 4324 6662 4380
rect 6598 4320 6662 4324
rect 1630 3836 1694 3840
rect 1630 3780 1634 3836
rect 1634 3780 1690 3836
rect 1690 3780 1694 3836
rect 1630 3776 1694 3780
rect 1710 3836 1774 3840
rect 1710 3780 1714 3836
rect 1714 3780 1770 3836
rect 1770 3780 1774 3836
rect 1710 3776 1774 3780
rect 1790 3836 1854 3840
rect 1790 3780 1794 3836
rect 1794 3780 1850 3836
rect 1850 3780 1854 3836
rect 1790 3776 1854 3780
rect 1870 3836 1934 3840
rect 1870 3780 1874 3836
rect 1874 3780 1930 3836
rect 1930 3780 1934 3836
rect 1870 3776 1934 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 3146 3836 3210 3840
rect 3146 3780 3150 3836
rect 3150 3780 3206 3836
rect 3206 3780 3210 3836
rect 3146 3776 3210 3780
rect 3226 3836 3290 3840
rect 3226 3780 3230 3836
rect 3230 3780 3286 3836
rect 3286 3780 3290 3836
rect 3226 3776 3290 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 4422 3836 4486 3840
rect 4422 3780 4426 3836
rect 4426 3780 4482 3836
rect 4482 3780 4486 3836
rect 4422 3776 4486 3780
rect 4502 3836 4566 3840
rect 4502 3780 4506 3836
rect 4506 3780 4562 3836
rect 4562 3780 4566 3836
rect 4502 3776 4566 3780
rect 4582 3836 4646 3840
rect 4582 3780 4586 3836
rect 4586 3780 4642 3836
rect 4642 3780 4646 3836
rect 4582 3776 4646 3780
rect 5698 3836 5762 3840
rect 5698 3780 5702 3836
rect 5702 3780 5758 3836
rect 5758 3780 5762 3836
rect 5698 3776 5762 3780
rect 5778 3836 5842 3840
rect 5778 3780 5782 3836
rect 5782 3780 5838 3836
rect 5838 3780 5842 3836
rect 5778 3776 5842 3780
rect 5858 3836 5922 3840
rect 5858 3780 5862 3836
rect 5862 3780 5918 3836
rect 5918 3780 5922 3836
rect 5858 3776 5922 3780
rect 5938 3836 6002 3840
rect 5938 3780 5942 3836
rect 5942 3780 5998 3836
rect 5998 3780 6002 3836
rect 5938 3776 6002 3780
rect 2290 3292 2354 3296
rect 2290 3236 2294 3292
rect 2294 3236 2350 3292
rect 2350 3236 2354 3292
rect 2290 3232 2354 3236
rect 2370 3292 2434 3296
rect 2370 3236 2374 3292
rect 2374 3236 2430 3292
rect 2430 3236 2434 3292
rect 2370 3232 2434 3236
rect 2450 3292 2514 3296
rect 2450 3236 2454 3292
rect 2454 3236 2510 3292
rect 2510 3236 2514 3292
rect 2450 3232 2514 3236
rect 2530 3292 2594 3296
rect 2530 3236 2534 3292
rect 2534 3236 2590 3292
rect 2590 3236 2594 3292
rect 2530 3232 2594 3236
rect 3646 3292 3710 3296
rect 3646 3236 3650 3292
rect 3650 3236 3706 3292
rect 3706 3236 3710 3292
rect 3646 3232 3710 3236
rect 3726 3292 3790 3296
rect 3726 3236 3730 3292
rect 3730 3236 3786 3292
rect 3786 3236 3790 3292
rect 3726 3232 3790 3236
rect 3806 3292 3870 3296
rect 3806 3236 3810 3292
rect 3810 3236 3866 3292
rect 3866 3236 3870 3292
rect 3806 3232 3870 3236
rect 3886 3292 3950 3296
rect 3886 3236 3890 3292
rect 3890 3236 3946 3292
rect 3946 3236 3950 3292
rect 3886 3232 3950 3236
rect 5002 3292 5066 3296
rect 5002 3236 5006 3292
rect 5006 3236 5062 3292
rect 5062 3236 5066 3292
rect 5002 3232 5066 3236
rect 5082 3292 5146 3296
rect 5082 3236 5086 3292
rect 5086 3236 5142 3292
rect 5142 3236 5146 3292
rect 5082 3232 5146 3236
rect 5162 3292 5226 3296
rect 5162 3236 5166 3292
rect 5166 3236 5222 3292
rect 5222 3236 5226 3292
rect 5162 3232 5226 3236
rect 5242 3292 5306 3296
rect 5242 3236 5246 3292
rect 5246 3236 5302 3292
rect 5302 3236 5306 3292
rect 5242 3232 5306 3236
rect 6358 3292 6422 3296
rect 6358 3236 6362 3292
rect 6362 3236 6418 3292
rect 6418 3236 6422 3292
rect 6358 3232 6422 3236
rect 6438 3292 6502 3296
rect 6438 3236 6442 3292
rect 6442 3236 6498 3292
rect 6498 3236 6502 3292
rect 6438 3232 6502 3236
rect 6518 3292 6582 3296
rect 6518 3236 6522 3292
rect 6522 3236 6578 3292
rect 6578 3236 6582 3292
rect 6518 3232 6582 3236
rect 6598 3292 6662 3296
rect 6598 3236 6602 3292
rect 6602 3236 6658 3292
rect 6658 3236 6662 3292
rect 6598 3232 6662 3236
rect 1630 2748 1694 2752
rect 1630 2692 1634 2748
rect 1634 2692 1690 2748
rect 1690 2692 1694 2748
rect 1630 2688 1694 2692
rect 1710 2748 1774 2752
rect 1710 2692 1714 2748
rect 1714 2692 1770 2748
rect 1770 2692 1774 2748
rect 1710 2688 1774 2692
rect 1790 2748 1854 2752
rect 1790 2692 1794 2748
rect 1794 2692 1850 2748
rect 1850 2692 1854 2748
rect 1790 2688 1854 2692
rect 1870 2748 1934 2752
rect 1870 2692 1874 2748
rect 1874 2692 1930 2748
rect 1930 2692 1934 2748
rect 1870 2688 1934 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 3146 2748 3210 2752
rect 3146 2692 3150 2748
rect 3150 2692 3206 2748
rect 3206 2692 3210 2748
rect 3146 2688 3210 2692
rect 3226 2748 3290 2752
rect 3226 2692 3230 2748
rect 3230 2692 3286 2748
rect 3286 2692 3290 2748
rect 3226 2688 3290 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 4422 2748 4486 2752
rect 4422 2692 4426 2748
rect 4426 2692 4482 2748
rect 4482 2692 4486 2748
rect 4422 2688 4486 2692
rect 4502 2748 4566 2752
rect 4502 2692 4506 2748
rect 4506 2692 4562 2748
rect 4562 2692 4566 2748
rect 4502 2688 4566 2692
rect 4582 2748 4646 2752
rect 4582 2692 4586 2748
rect 4586 2692 4642 2748
rect 4642 2692 4646 2748
rect 4582 2688 4646 2692
rect 5698 2748 5762 2752
rect 5698 2692 5702 2748
rect 5702 2692 5758 2748
rect 5758 2692 5762 2748
rect 5698 2688 5762 2692
rect 5778 2748 5842 2752
rect 5778 2692 5782 2748
rect 5782 2692 5838 2748
rect 5838 2692 5842 2748
rect 5778 2688 5842 2692
rect 5858 2748 5922 2752
rect 5858 2692 5862 2748
rect 5862 2692 5918 2748
rect 5918 2692 5922 2748
rect 5858 2688 5922 2692
rect 5938 2748 6002 2752
rect 5938 2692 5942 2748
rect 5942 2692 5998 2748
rect 5998 2692 6002 2748
rect 5938 2688 6002 2692
rect 2290 2204 2354 2208
rect 2290 2148 2294 2204
rect 2294 2148 2350 2204
rect 2350 2148 2354 2204
rect 2290 2144 2354 2148
rect 2370 2204 2434 2208
rect 2370 2148 2374 2204
rect 2374 2148 2430 2204
rect 2430 2148 2434 2204
rect 2370 2144 2434 2148
rect 2450 2204 2514 2208
rect 2450 2148 2454 2204
rect 2454 2148 2510 2204
rect 2510 2148 2514 2204
rect 2450 2144 2514 2148
rect 2530 2204 2594 2208
rect 2530 2148 2534 2204
rect 2534 2148 2590 2204
rect 2590 2148 2594 2204
rect 2530 2144 2594 2148
rect 3646 2204 3710 2208
rect 3646 2148 3650 2204
rect 3650 2148 3706 2204
rect 3706 2148 3710 2204
rect 3646 2144 3710 2148
rect 3726 2204 3790 2208
rect 3726 2148 3730 2204
rect 3730 2148 3786 2204
rect 3786 2148 3790 2204
rect 3726 2144 3790 2148
rect 3806 2204 3870 2208
rect 3806 2148 3810 2204
rect 3810 2148 3866 2204
rect 3866 2148 3870 2204
rect 3806 2144 3870 2148
rect 3886 2204 3950 2208
rect 3886 2148 3890 2204
rect 3890 2148 3946 2204
rect 3946 2148 3950 2204
rect 3886 2144 3950 2148
rect 5002 2204 5066 2208
rect 5002 2148 5006 2204
rect 5006 2148 5062 2204
rect 5062 2148 5066 2204
rect 5002 2144 5066 2148
rect 5082 2204 5146 2208
rect 5082 2148 5086 2204
rect 5086 2148 5142 2204
rect 5142 2148 5146 2204
rect 5082 2144 5146 2148
rect 5162 2204 5226 2208
rect 5162 2148 5166 2204
rect 5166 2148 5222 2204
rect 5222 2148 5226 2204
rect 5162 2144 5226 2148
rect 5242 2204 5306 2208
rect 5242 2148 5246 2204
rect 5246 2148 5302 2204
rect 5302 2148 5306 2204
rect 5242 2144 5306 2148
rect 6358 2204 6422 2208
rect 6358 2148 6362 2204
rect 6362 2148 6418 2204
rect 6418 2148 6422 2204
rect 6358 2144 6422 2148
rect 6438 2204 6502 2208
rect 6438 2148 6442 2204
rect 6442 2148 6498 2204
rect 6498 2148 6502 2204
rect 6438 2144 6502 2148
rect 6518 2204 6582 2208
rect 6518 2148 6522 2204
rect 6522 2148 6578 2204
rect 6578 2148 6582 2204
rect 6518 2144 6582 2148
rect 6598 2204 6662 2208
rect 6598 2148 6602 2204
rect 6602 2148 6658 2204
rect 6658 2148 6662 2204
rect 6598 2144 6662 2148
<< metal4 >>
rect 2282 7710 2602 7752
rect 1622 7104 1942 7664
rect 1622 7040 1630 7104
rect 1694 7050 1710 7104
rect 1774 7050 1790 7104
rect 1854 7050 1870 7104
rect 1934 7040 1942 7104
rect 1622 6814 1664 7040
rect 1900 6814 1942 7040
rect 1622 6016 1942 6814
rect 1622 5952 1630 6016
rect 1694 5952 1710 6016
rect 1774 5952 1790 6016
rect 1854 5952 1870 6016
rect 1934 5952 1942 6016
rect 1622 5691 1942 5952
rect 1622 5455 1664 5691
rect 1900 5455 1942 5691
rect 1622 4928 1942 5455
rect 1622 4864 1630 4928
rect 1694 4864 1710 4928
rect 1774 4864 1790 4928
rect 1854 4864 1870 4928
rect 1934 4864 1942 4928
rect 1622 4332 1942 4864
rect 1622 4096 1664 4332
rect 1900 4096 1942 4332
rect 1622 3840 1942 4096
rect 1622 3776 1630 3840
rect 1694 3776 1710 3840
rect 1774 3776 1790 3840
rect 1854 3776 1870 3840
rect 1934 3776 1942 3840
rect 1622 2973 1942 3776
rect 1622 2752 1664 2973
rect 1900 2752 1942 2973
rect 1622 2688 1630 2752
rect 1694 2688 1710 2737
rect 1774 2688 1790 2737
rect 1854 2688 1870 2737
rect 1934 2688 1942 2752
rect 1622 2128 1942 2688
rect 2282 7648 2324 7710
rect 2560 7648 2602 7710
rect 3638 7710 3958 7752
rect 2282 7584 2290 7648
rect 2594 7584 2602 7648
rect 2282 7474 2324 7584
rect 2560 7474 2602 7584
rect 2282 6560 2602 7474
rect 2282 6496 2290 6560
rect 2354 6496 2370 6560
rect 2434 6496 2450 6560
rect 2514 6496 2530 6560
rect 2594 6496 2602 6560
rect 2282 6351 2602 6496
rect 2282 6115 2324 6351
rect 2560 6115 2602 6351
rect 2282 5472 2602 6115
rect 2282 5408 2290 5472
rect 2354 5408 2370 5472
rect 2434 5408 2450 5472
rect 2514 5408 2530 5472
rect 2594 5408 2602 5472
rect 2282 4992 2602 5408
rect 2282 4756 2324 4992
rect 2560 4756 2602 4992
rect 2282 4384 2602 4756
rect 2282 4320 2290 4384
rect 2354 4320 2370 4384
rect 2434 4320 2450 4384
rect 2514 4320 2530 4384
rect 2594 4320 2602 4384
rect 2282 3633 2602 4320
rect 2282 3397 2324 3633
rect 2560 3397 2602 3633
rect 2282 3296 2602 3397
rect 2282 3232 2290 3296
rect 2354 3232 2370 3296
rect 2434 3232 2450 3296
rect 2514 3232 2530 3296
rect 2594 3232 2602 3296
rect 2282 2208 2602 3232
rect 2282 2144 2290 2208
rect 2354 2144 2370 2208
rect 2434 2144 2450 2208
rect 2514 2144 2530 2208
rect 2594 2144 2602 2208
rect 2282 2128 2602 2144
rect 2978 7104 3298 7664
rect 2978 7040 2986 7104
rect 3050 7050 3066 7104
rect 3130 7050 3146 7104
rect 3210 7050 3226 7104
rect 3290 7040 3298 7104
rect 2978 6814 3020 7040
rect 3256 6814 3298 7040
rect 2978 6016 3298 6814
rect 2978 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3146 6016
rect 3210 5952 3226 6016
rect 3290 5952 3298 6016
rect 2978 5691 3298 5952
rect 2978 5455 3020 5691
rect 3256 5455 3298 5691
rect 2978 4928 3298 5455
rect 2978 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3146 4928
rect 3210 4864 3226 4928
rect 3290 4864 3298 4928
rect 2978 4332 3298 4864
rect 2978 4096 3020 4332
rect 3256 4096 3298 4332
rect 2978 3840 3298 4096
rect 2978 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3146 3840
rect 3210 3776 3226 3840
rect 3290 3776 3298 3840
rect 2978 2973 3298 3776
rect 2978 2752 3020 2973
rect 3256 2752 3298 2973
rect 2978 2688 2986 2752
rect 3050 2688 3066 2737
rect 3130 2688 3146 2737
rect 3210 2688 3226 2737
rect 3290 2688 3298 2752
rect 2978 2128 3298 2688
rect 3638 7648 3680 7710
rect 3916 7648 3958 7710
rect 4994 7710 5314 7752
rect 3638 7584 3646 7648
rect 3950 7584 3958 7648
rect 3638 7474 3680 7584
rect 3916 7474 3958 7584
rect 3638 6560 3958 7474
rect 3638 6496 3646 6560
rect 3710 6496 3726 6560
rect 3790 6496 3806 6560
rect 3870 6496 3886 6560
rect 3950 6496 3958 6560
rect 3638 6351 3958 6496
rect 3638 6115 3680 6351
rect 3916 6115 3958 6351
rect 3638 5472 3958 6115
rect 3638 5408 3646 5472
rect 3710 5408 3726 5472
rect 3790 5408 3806 5472
rect 3870 5408 3886 5472
rect 3950 5408 3958 5472
rect 3638 4992 3958 5408
rect 3638 4756 3680 4992
rect 3916 4756 3958 4992
rect 3638 4384 3958 4756
rect 3638 4320 3646 4384
rect 3710 4320 3726 4384
rect 3790 4320 3806 4384
rect 3870 4320 3886 4384
rect 3950 4320 3958 4384
rect 3638 3633 3958 4320
rect 3638 3397 3680 3633
rect 3916 3397 3958 3633
rect 3638 3296 3958 3397
rect 3638 3232 3646 3296
rect 3710 3232 3726 3296
rect 3790 3232 3806 3296
rect 3870 3232 3886 3296
rect 3950 3232 3958 3296
rect 3638 2208 3958 3232
rect 3638 2144 3646 2208
rect 3710 2144 3726 2208
rect 3790 2144 3806 2208
rect 3870 2144 3886 2208
rect 3950 2144 3958 2208
rect 3638 2128 3958 2144
rect 4334 7104 4654 7664
rect 4334 7040 4342 7104
rect 4406 7050 4422 7104
rect 4486 7050 4502 7104
rect 4566 7050 4582 7104
rect 4646 7040 4654 7104
rect 4334 6814 4376 7040
rect 4612 6814 4654 7040
rect 4334 6016 4654 6814
rect 4334 5952 4342 6016
rect 4406 5952 4422 6016
rect 4486 5952 4502 6016
rect 4566 5952 4582 6016
rect 4646 5952 4654 6016
rect 4334 5691 4654 5952
rect 4334 5455 4376 5691
rect 4612 5455 4654 5691
rect 4334 4928 4654 5455
rect 4334 4864 4342 4928
rect 4406 4864 4422 4928
rect 4486 4864 4502 4928
rect 4566 4864 4582 4928
rect 4646 4864 4654 4928
rect 4334 4332 4654 4864
rect 4334 4096 4376 4332
rect 4612 4096 4654 4332
rect 4334 3840 4654 4096
rect 4334 3776 4342 3840
rect 4406 3776 4422 3840
rect 4486 3776 4502 3840
rect 4566 3776 4582 3840
rect 4646 3776 4654 3840
rect 4334 2973 4654 3776
rect 4334 2752 4376 2973
rect 4612 2752 4654 2973
rect 4334 2688 4342 2752
rect 4406 2688 4422 2737
rect 4486 2688 4502 2737
rect 4566 2688 4582 2737
rect 4646 2688 4654 2752
rect 4334 2128 4654 2688
rect 4994 7648 5036 7710
rect 5272 7648 5314 7710
rect 6350 7710 6670 7752
rect 4994 7584 5002 7648
rect 5306 7584 5314 7648
rect 4994 7474 5036 7584
rect 5272 7474 5314 7584
rect 4994 6560 5314 7474
rect 4994 6496 5002 6560
rect 5066 6496 5082 6560
rect 5146 6496 5162 6560
rect 5226 6496 5242 6560
rect 5306 6496 5314 6560
rect 4994 6351 5314 6496
rect 4994 6115 5036 6351
rect 5272 6115 5314 6351
rect 4994 5472 5314 6115
rect 4994 5408 5002 5472
rect 5066 5408 5082 5472
rect 5146 5408 5162 5472
rect 5226 5408 5242 5472
rect 5306 5408 5314 5472
rect 4994 4992 5314 5408
rect 4994 4756 5036 4992
rect 5272 4756 5314 4992
rect 4994 4384 5314 4756
rect 4994 4320 5002 4384
rect 5066 4320 5082 4384
rect 5146 4320 5162 4384
rect 5226 4320 5242 4384
rect 5306 4320 5314 4384
rect 4994 3633 5314 4320
rect 4994 3397 5036 3633
rect 5272 3397 5314 3633
rect 4994 3296 5314 3397
rect 4994 3232 5002 3296
rect 5066 3232 5082 3296
rect 5146 3232 5162 3296
rect 5226 3232 5242 3296
rect 5306 3232 5314 3296
rect 4994 2208 5314 3232
rect 4994 2144 5002 2208
rect 5066 2144 5082 2208
rect 5146 2144 5162 2208
rect 5226 2144 5242 2208
rect 5306 2144 5314 2208
rect 4994 2128 5314 2144
rect 5690 7104 6010 7664
rect 5690 7040 5698 7104
rect 5762 7050 5778 7104
rect 5842 7050 5858 7104
rect 5922 7050 5938 7104
rect 6002 7040 6010 7104
rect 5690 6814 5732 7040
rect 5968 6814 6010 7040
rect 5690 6016 6010 6814
rect 5690 5952 5698 6016
rect 5762 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5938 6016
rect 6002 5952 6010 6016
rect 5690 5691 6010 5952
rect 5690 5455 5732 5691
rect 5968 5455 6010 5691
rect 5690 4928 6010 5455
rect 5690 4864 5698 4928
rect 5762 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5938 4928
rect 6002 4864 6010 4928
rect 5690 4332 6010 4864
rect 5690 4096 5732 4332
rect 5968 4096 6010 4332
rect 5690 3840 6010 4096
rect 5690 3776 5698 3840
rect 5762 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5938 3840
rect 6002 3776 6010 3840
rect 5690 2973 6010 3776
rect 5690 2752 5732 2973
rect 5968 2752 6010 2973
rect 5690 2688 5698 2752
rect 5762 2688 5778 2737
rect 5842 2688 5858 2737
rect 5922 2688 5938 2737
rect 6002 2688 6010 2752
rect 5690 2128 6010 2688
rect 6350 7648 6392 7710
rect 6628 7648 6670 7710
rect 6350 7584 6358 7648
rect 6662 7584 6670 7648
rect 6350 7474 6392 7584
rect 6628 7474 6670 7584
rect 6350 6560 6670 7474
rect 6350 6496 6358 6560
rect 6422 6496 6438 6560
rect 6502 6496 6518 6560
rect 6582 6496 6598 6560
rect 6662 6496 6670 6560
rect 6350 6351 6670 6496
rect 6350 6115 6392 6351
rect 6628 6115 6670 6351
rect 6350 5472 6670 6115
rect 6350 5408 6358 5472
rect 6422 5408 6438 5472
rect 6502 5408 6518 5472
rect 6582 5408 6598 5472
rect 6662 5408 6670 5472
rect 6350 4992 6670 5408
rect 6350 4756 6392 4992
rect 6628 4756 6670 4992
rect 6350 4384 6670 4756
rect 6350 4320 6358 4384
rect 6422 4320 6438 4384
rect 6502 4320 6518 4384
rect 6582 4320 6598 4384
rect 6662 4320 6670 4384
rect 6350 3633 6670 4320
rect 6350 3397 6392 3633
rect 6628 3397 6670 3633
rect 6350 3296 6670 3397
rect 6350 3232 6358 3296
rect 6422 3232 6438 3296
rect 6502 3232 6518 3296
rect 6582 3232 6598 3296
rect 6662 3232 6670 3296
rect 6350 2208 6670 3232
rect 6350 2144 6358 2208
rect 6422 2144 6438 2208
rect 6502 2144 6518 2208
rect 6582 2144 6598 2208
rect 6662 2144 6670 2208
rect 6350 2128 6670 2144
<< via4 >>
rect 1664 7040 1694 7050
rect 1694 7040 1710 7050
rect 1710 7040 1774 7050
rect 1774 7040 1790 7050
rect 1790 7040 1854 7050
rect 1854 7040 1870 7050
rect 1870 7040 1900 7050
rect 1664 6814 1900 7040
rect 1664 5455 1900 5691
rect 1664 4096 1900 4332
rect 1664 2752 1900 2973
rect 1664 2737 1694 2752
rect 1694 2737 1710 2752
rect 1710 2737 1774 2752
rect 1774 2737 1790 2752
rect 1790 2737 1854 2752
rect 1854 2737 1870 2752
rect 1870 2737 1900 2752
rect 2324 7648 2560 7710
rect 2324 7584 2354 7648
rect 2354 7584 2370 7648
rect 2370 7584 2434 7648
rect 2434 7584 2450 7648
rect 2450 7584 2514 7648
rect 2514 7584 2530 7648
rect 2530 7584 2560 7648
rect 2324 7474 2560 7584
rect 2324 6115 2560 6351
rect 2324 4756 2560 4992
rect 2324 3397 2560 3633
rect 3020 7040 3050 7050
rect 3050 7040 3066 7050
rect 3066 7040 3130 7050
rect 3130 7040 3146 7050
rect 3146 7040 3210 7050
rect 3210 7040 3226 7050
rect 3226 7040 3256 7050
rect 3020 6814 3256 7040
rect 3020 5455 3256 5691
rect 3020 4096 3256 4332
rect 3020 2752 3256 2973
rect 3020 2737 3050 2752
rect 3050 2737 3066 2752
rect 3066 2737 3130 2752
rect 3130 2737 3146 2752
rect 3146 2737 3210 2752
rect 3210 2737 3226 2752
rect 3226 2737 3256 2752
rect 3680 7648 3916 7710
rect 3680 7584 3710 7648
rect 3710 7584 3726 7648
rect 3726 7584 3790 7648
rect 3790 7584 3806 7648
rect 3806 7584 3870 7648
rect 3870 7584 3886 7648
rect 3886 7584 3916 7648
rect 3680 7474 3916 7584
rect 3680 6115 3916 6351
rect 3680 4756 3916 4992
rect 3680 3397 3916 3633
rect 4376 7040 4406 7050
rect 4406 7040 4422 7050
rect 4422 7040 4486 7050
rect 4486 7040 4502 7050
rect 4502 7040 4566 7050
rect 4566 7040 4582 7050
rect 4582 7040 4612 7050
rect 4376 6814 4612 7040
rect 4376 5455 4612 5691
rect 4376 4096 4612 4332
rect 4376 2752 4612 2973
rect 4376 2737 4406 2752
rect 4406 2737 4422 2752
rect 4422 2737 4486 2752
rect 4486 2737 4502 2752
rect 4502 2737 4566 2752
rect 4566 2737 4582 2752
rect 4582 2737 4612 2752
rect 5036 7648 5272 7710
rect 5036 7584 5066 7648
rect 5066 7584 5082 7648
rect 5082 7584 5146 7648
rect 5146 7584 5162 7648
rect 5162 7584 5226 7648
rect 5226 7584 5242 7648
rect 5242 7584 5272 7648
rect 5036 7474 5272 7584
rect 5036 6115 5272 6351
rect 5036 4756 5272 4992
rect 5036 3397 5272 3633
rect 5732 7040 5762 7050
rect 5762 7040 5778 7050
rect 5778 7040 5842 7050
rect 5842 7040 5858 7050
rect 5858 7040 5922 7050
rect 5922 7040 5938 7050
rect 5938 7040 5968 7050
rect 5732 6814 5968 7040
rect 5732 5455 5968 5691
rect 5732 4096 5968 4332
rect 5732 2752 5968 2973
rect 5732 2737 5762 2752
rect 5762 2737 5778 2752
rect 5778 2737 5842 2752
rect 5842 2737 5858 2752
rect 5858 2737 5922 2752
rect 5922 2737 5938 2752
rect 5938 2737 5968 2752
rect 6392 7648 6628 7710
rect 6392 7584 6422 7648
rect 6422 7584 6438 7648
rect 6438 7584 6502 7648
rect 6502 7584 6518 7648
rect 6518 7584 6582 7648
rect 6582 7584 6598 7648
rect 6598 7584 6628 7648
rect 6392 7474 6628 7584
rect 6392 6115 6628 6351
rect 6392 4756 6628 4992
rect 6392 3397 6628 3633
<< metal5 >>
rect 1056 7710 6670 7752
rect 1056 7474 2324 7710
rect 2560 7474 3680 7710
rect 3916 7474 5036 7710
rect 5272 7474 6392 7710
rect 6628 7474 6670 7710
rect 1056 7432 6670 7474
rect 1056 7050 6580 7092
rect 1056 6814 1664 7050
rect 1900 6814 3020 7050
rect 3256 6814 4376 7050
rect 4612 6814 5732 7050
rect 5968 6814 6580 7050
rect 1056 6772 6580 6814
rect 1056 6351 6670 6393
rect 1056 6115 2324 6351
rect 2560 6115 3680 6351
rect 3916 6115 5036 6351
rect 5272 6115 6392 6351
rect 6628 6115 6670 6351
rect 1056 6073 6670 6115
rect 1056 5691 6580 5733
rect 1056 5455 1664 5691
rect 1900 5455 3020 5691
rect 3256 5455 4376 5691
rect 4612 5455 5732 5691
rect 5968 5455 6580 5691
rect 1056 5413 6580 5455
rect 1056 4992 6670 5034
rect 1056 4756 2324 4992
rect 2560 4756 3680 4992
rect 3916 4756 5036 4992
rect 5272 4756 6392 4992
rect 6628 4756 6670 4992
rect 1056 4714 6670 4756
rect 1056 4332 6580 4374
rect 1056 4096 1664 4332
rect 1900 4096 3020 4332
rect 3256 4096 4376 4332
rect 4612 4096 5732 4332
rect 5968 4096 6580 4332
rect 1056 4054 6580 4096
rect 1056 3633 6670 3675
rect 1056 3397 2324 3633
rect 2560 3397 3680 3633
rect 3916 3397 5036 3633
rect 5272 3397 6392 3633
rect 6628 3397 6670 3633
rect 1056 3355 6670 3397
rect 1056 2973 6580 3015
rect 1056 2737 1664 2973
rect 1900 2737 3020 2973
rect 3256 2737 4376 2973
rect 4612 2737 5732 2973
rect 5968 2737 6580 2973
rect 1056 2695 6580 2737
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_29
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_41
timestamp 0
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 0
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pes_sipo_1
timestamp 0
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pes_sipo_2
timestamp 0
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pes_sipo_3
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pes_sipo_4
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_21
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_22
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_23
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_24
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_25
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
<< labels >>
rlabel metal2 s 3887 7616 3887 7616 4 VGND
rlabel metal1 s 3818 7072 3818 7072 4 VPWR
rlabel metal3 s 6210 6171 6210 6171 4 net1
rlabel metal2 s 6210 4913 6210 4913 4 net2
rlabel metal2 s 6210 4369 6210 4369 4 net3
rlabel metal1 s 6486 5678 6486 5678 4 net4
flabel metal5 s 1056 7432 6670 7752 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6073 6670 6393 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4714 6670 5034 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3355 6670 3675 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 6350 2128 6670 7752 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4994 2128 5314 7752 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3638 2128 3958 7752 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2282 2128 2602 7752 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6772 6580 7092 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5413 6580 5733 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4054 6580 4374 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 2695 6580 3015 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 5690 2128 6010 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4334 2128 4654 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2978 2128 3298 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1622 2128 1942 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 b
port 3 nsew
flabel metal2 s 662 0 718 800 0 FreeSans 280 90 0 0 clk
port 4 nsew
flabel metal3 s 6888 6128 7688 6248 0 FreeSans 600 0 0 0 q[0]
port 5 nsew
flabel metal3 s 6888 4768 7688 4888 0 FreeSans 600 0 0 0 q[1]
port 6 nsew
flabel metal3 s 6888 4088 7688 4208 0 FreeSans 600 0 0 0 q[2]
port 7 nsew
flabel metal3 s 6888 5448 7688 5568 0 FreeSans 600 0 0 0 q[3]
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 7688 9832
<< end >>
